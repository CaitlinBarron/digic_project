
-- 
-- Definition of  MAC
-- 
--      Sun Dec  8 19:15:39 2019
--      
--      LeonardoSpectrum Level 3, 2008b.3
-- 

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity Multiplier_32 is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      Product : OUT std_logic_vector (31 DOWNTO 0)) ;
end Multiplier_32 ;

architecture structural of Multiplier_32 is
   signal Product_0_EXMPLR, nx14, nx20, nx36, nx44, nx52, nx68, nx70, nx74, 
      nx88, nx96, nx112, nx114, nx122, nx128, nx144, nx152, nx168, nx170, 
      nx180, nx188, nx196, nx212, nx220, nx236, nx238, nx248, nx250, nx254, 
      nx268, nx276, nx292, nx300, nx316, nx318, nx328, nx330, nx338, nx344, 
      nx360, nx368, nx384, nx392, nx408, nx410, nx420, nx422, nx432, nx440, 
      nx448, nx464, nx472, nx488, nx496, nx512, nx514, nx524, nx526, nx536, 
      nx538, nx542, nx556, nx564, nx580, nx588, nx604, nx612, nx628, nx630, 
      nx640, nx642, nx652, nx654, nx662, nx668, nx684, nx692, nx708, nx716, 
      nx732, nx740, nx756, nx758, nx768, nx770, nx780, nx782, nx792, nx800, 
      nx808, nx824, nx832, nx848, nx856, nx872, nx880, nx896, nx898, nx908, 
      nx910, nx920, nx922, nx932, nx934, nx938, nx952, nx960, nx976, nx984, 
      nx1000, nx1008, nx1024, nx1032, nx1048, nx1050, nx1060, nx1062, nx1072, 
      nx1074, nx1084, nx1086, nx1094, nx1100, nx1116, nx1124, nx1140, nx1148, 
      nx1164, nx1172, nx1188, nx1196, nx1212, nx1214, nx1224, nx1226, nx1236, 
      nx1238, nx1248, nx1250, nx1260, nx1262, nx1268, nx1274, nx1290, nx1298, 
      nx1314, nx1322, nx1338, nx1346, nx1362, nx1370, nx1382, nx1390, nx1392, 
      nx1402, nx1404, nx1414, nx1416, nx1426, nx1428, nx1438, nx1440, nx1446, 
      nx1452, nx1458, nx1466, nx1474, nx1482, nx1490, nx1498, nx1506, nx1514, 
      nx1522, nx1530, nx1538, nx1546, nx1558, nx1560, nx1562, nx1564, nx1570, 
      nx1572, nx1574, nx1576, nx1582, nx1584, nx1586, nx1588, nx1594, nx1596, 
      nx1598, nx1600, nx1602, nx1604, nx1622, nx1630, nx1654, nx1662, nx1670, 
      nx1678, nx1702, nx1710, nx1718, nx1720, nx1734, nx1736, nx1738, nx1740, 
      nx1742, nx1744, nx1758, nx1760, nx1762, nx1764, nx1770, nx1776, nx1782, 
      nx1790, nx1798, nx1830, nx1838, nx1846, nx1854, nx1862, nx1870, nx1872, 
      nx1874, nx1876, nx1882, nx1884, nx1902, nx1904, nx1910, nx1912, nx1924, 
      nx1938, nx1946, nx1954, nx1962, nx1978, nx1986, nx1994, nx2002, nx2010, 
      nx2012, nx2014, nx2016, nx2018, nx2020, nx2030, nx2032, nx2038, nx2040, 
      nx2048, nx2054, nx2060, nx2074, nx2082, nx2090, nx2098, nx2106, nx2114, 
      nx2122, nx2130, nx2138, nx2140, nx2142, nx2144, nx2146, nx2148, nx2150, 
      nx2152, nx2158, nx2160, nx2162, nx2164, nx2170, nx2172, nx2184, nx2206, 
      nx2214, nx2222, nx2230, nx2238, nx2246, nx2254, nx2256, nx2258, nx2260, 
      nx2262, nx2264, nx2266, nx2268, nx2270, nx2272, nx2284, nx2290, nx2296, 
      nx2302, nx2310, nx2318, nx2326, nx2334, nx2342, nx2350, nx2358, nx2360, 
      nx2362, nx2364, nx2366, nx2368, nx2370, nx2372, nx2374, nx2376, nx2378, 
      nx2380, nx2382, nx2384, nx2402, nx2410, nx2418, nx2426, nx2434, nx2442, 
      nx2450, nx2452, nx2454, nx2456, nx2458, nx2460, nx2462, nx2464, nx2466, 
      nx2468, nx2470, nx2472, nx2478, nx2484, nx2490, nx2498, nx2506, nx2514, 
      nx2522, nx2530, nx2532, nx2534, nx2536, nx2538, nx2540, nx2542, nx2544, 
      nx2546, nx2548, nx2566, nx2574, nx2582, nx2590, nx2598, nx2600, nx2602, 
      nx2604, nx2606, nx2608, nx2610, nx2612, nx2618, nx2624, nx2630, nx2638, 
      nx2646, nx2654, nx2656, nx2658, nx2660, nx2662, nx2664, nx2682, nx2690, 
      nx2698, nx2700, nx2702, nx2704, nx2710, nx2716, nx2722, nx2730, nx2732, 
      nx2738, nx2744, nx2748, nx1551, nx1553, nx1559, nx1561, nx1563, nx1567, 
      nx1569, nx1571, nx1573, nx1579, nx1581, nx1583, nx1587, nx1589, nx1591, 
      nx1593, nx1595, nx1597, nx1599, nx1601, nx1605, nx1607, nx1611, nx1613, 
      nx1615, nx1617, nx1621, nx1627, nx1629, nx1631, nx1633, nx1635, nx1637, 
      nx1639, nx1641, nx1643, nx1645, nx1647, nx1653, nx1657, nx1659, nx1661, 
      nx1667, nx1669, nx1671, nx1673, nx1677, nx1679, nx1681, nx1683, nx1685, 
      nx1687, nx1689, nx1691, nx1693, nx1695, nx1699, nx1703, nx1709, nx1715, 
      nx1717, nx1719, nx1721, nx1723, nx1725, nx1727, nx1731, nx1733, nx1735, 
      nx1737, nx1741, nx1743, nx1749, nx1753, nx1755, nx1757, nx1763, nx1765, 
      nx1767, nx1769, nx1773, nx1775, nx1777, nx1779, nx1781, nx1785, nx1787, 
      nx1789, nx1791, nx1795, nx1799, nx1805, nx1807, nx1809, nx1811, nx1813, 
      nx1815, nx1817, nx1821, nx1825, nx1831, nx1837, nx1839, nx1841, nx1843, 
      nx1845, nx1847, nx1849, nx1851, nx1855, nx1857, nx1859, nx1865, nx1867, 
      nx1871, nx1873, nx1879, nx1883, nx1885, nx1887, nx1893, nx1895, nx1897, 
      nx1899, nx1903, nx1905, nx1907, nx1909, nx1911, nx1915, nx1917, nx1919, 
      nx1921, nx1923, nx1927, nx1933, nx1935, nx1937, nx1939, nx1941, nx1943, 
      nx1945, nx1949, nx1953, nx1959, nx1961, nx1963, nx1965, nx1967, nx1969, 
      nx1971, nx1975, nx1979, nx1985, nx1991, nx1993, nx1995, nx1997, nx1999, 
      nx2001, nx2003, nx2005, nx2011, nx2013, nx2017, nx2019, nx2025, nx2027, 
      nx2031, nx2033, nx2039, nx2043, nx2045, nx2047, nx2053, nx2055, nx2057, 
      nx2059, nx2063, nx2065, nx2067, nx2069, nx2071, nx2075, nx2077, nx2079, 
      nx2081, nx2083, nx2087, nx2089, nx2091, nx2093, nx2095, nx2097, nx2099, 
      nx2101, nx2103, nx2105, nx2109, nx2113, nx2119, nx2121, nx2123, nx2125, 
      nx2127, nx2129, nx2131, nx2135, nx2139, nx2145, nx2147, nx2149, nx2151, 
      nx2153, nx2155, nx2157, nx2161, nx2165, nx2171, nx2177, nx2179, nx2181, 
      nx2183, nx2185, nx2187, nx2189, nx2193, nx2195, nx2197, nx2199, nx2203, 
      nx2205, nx2211, nx2213, nx2217, nx2219, nx2225, nx2227, nx2231, nx2233, 
      nx2239, nx2243, nx2245, nx2247, nx2253, nx2255, nx2257, nx2259, nx2263, 
      nx2265, nx2267, nx2269, nx2271, nx2275, nx2277, nx2279, nx2281, nx2283, 
      nx2287, nx2289, nx2291, nx2293, nx2295, nx2299, nx2301, nx2303, nx2305, 
      nx2309, nx2313, nx2319, nx2321, nx2323, nx2325, nx2327, nx2329, nx2331, 
      nx2335, nx2339, nx2345, nx2347, nx2349, nx2351, nx2353, nx2355, nx2357, 
      nx2361, nx2365, nx2371, nx2373, nx2375, nx2377, nx2379, nx2381, nx2383, 
      nx2387, nx2391, nx2397, nx2403, nx2405, nx2407, nx2409, nx2411, nx2413, 
      nx2415, nx2419, nx2423, nx2427, nx2431, nx2435, nx2439, nx2443, nx2447, 
      nx2451, nx2453, nx2455, nx2461, nx2465, nx2469, nx2473, nx2479, nx2481, 
      nx2483, nx2485, nx2487, nx2489, nx2491, nx2493, nx2497, nx2501, nx2507, 
      nx2509, nx2511, nx2513, nx2515, nx2517, nx2519, nx2523, nx2527, nx2533, 
      nx2535, nx2537, nx2539, nx2541, nx2543, nx2545, nx2549, nx2553, nx2559, 
      nx2561, nx2563, nx2565, nx2567, nx2569, nx2571, nx2575, nx2579, nx2585, 
      nx2591, nx2593, nx2595, nx2597, nx2599, nx2601, nx2603, nx2607, nx2637, 
      nx2639, nx2643, nx2645, nx2651, nx2653, nx2655, nx2657, nx2659, nx2661, 
      nx2663, nx2667, nx2671, nx2677, nx2679, nx2681, nx2683, nx2685, nx2687, 
      nx2689, nx2693, nx2697, nx2703, nx2705, nx2707, nx2709, nx2711, nx2713, 
      nx2715, nx2719, nx2723, nx2729, nx2731, nx2733, nx2735, nx2737, nx2739, 
      nx2741, nx2745, nx2749, nx2755, nx2761, nx2763, nx2765, nx2767, nx2769, 
      nx2775, nx2785, nx2787, nx2793, nx2797, nx2801, nx2807, nx2809, nx2811, 
      nx2813, nx2819, nx2823, nx2827, nx2833, nx2835, nx2837, nx2839, nx2845, 
      nx2849, nx2853, nx2859, nx2861, nx2863, nx2865, nx2871, nx2875, nx2879, 
      nx2883, nx2887, nx2889, nx2891, nx2893, nx2895, nx2897, nx2900, nx2907, 
      nx2910, nx2914, nx2918, nx2920, nx2924, nx2926, nx2928, nx2930, nx2932, 
      nx2934, nx2936, nx2938, nx2941, nx2943, nx2945, nx2948, nx2950, nx2955, 
      nx2958, nx2961, nx2964, nx2968, nx2972, nx2974, nx2978, nx2980, nx2982, 
      nx2984, nx2986, nx2988, nx2990, nx2992, nx2995, nx2997, nx2999, nx3002, 
      nx3004, nx3007, nx3011, nx3015, nx3017, nx3019, nx3023, nx3025, nx3028, 
      nx3033, nx3037, nx3039, nx3041, nx3045, nx3049, nx3051, nx3053, nx3055, 
      nx3057, nx3059, nx3061, nx3063, nx3066, nx3068, nx3070, nx3072, nx3075, 
      nx3077, nx3079, nx3082, nx3087, nx3091, nx3093, nx3095, nx3099, nx3102, 
      nx3105, nx3109, nx3111, nx3113, nx3115, nx3118, nx3123, nx3127, nx3129, 
      nx3131, nx3133, nx3135, nx3138, nx3141, nx3145, nx3147, nx3149, nx3153, 
      nx3157, nx3159, nx3161, nx3163, nx3165, nx3167, nx3169, nx3172, nx3175, 
      nx3178, nx3181, nx3184, nx3188, nx3192, nx3196, nx3198, nx3200, nx3204, 
      nx3206, nx3212, nx3214, nx3216, nx3218, nx3220, nx3223, nx3226, nx3229, 
      nx3232, nx3236, nx3238, nx3240, nx3242, nx3246, nx3249, nx3252, nx3255, 
      nx3259, nx3262, nx3266, nx3270, nx3274, nx3276, nx3278, nx3281, nx3286, 
      nx3288, nx3290, nx3292, nx3294, nx3296, nx3299, nx3301, nx3303, nx3306, 
      nx3311, nx3314, nx3317, nx3320, nx3324, nx3327, nx3331, nx3334, nx3338, 
      nx3342, nx3346, nx3348, nx3350, nx3354, nx3356, nx3360, nx3364, nx3367, 
      nx3370, nx3373, nx3377, nx3380, nx3384, nx3387, nx3391, nx3394, nx3398, 
      nx3402, nx3406, nx3408, nx3410, nx3413, nx3417, nx3420, nx3424, nx3427, 
      nx3431, nx3434, nx3438, nx3441, nx3445, nx3448, nx3452, nx3456, nx3460, 
      nx3462, nx3464, nx3468, nx3470, nx3473, nx3477, nx3481, nx3484, nx3488, 
      nx3491, nx3495, nx3498, nx3502, nx3506, nx3510, nx3512, nx3514, nx3517, 
      nx3521, nx3525, nx3529, nx3532, nx3536, nx3539, nx3543, nx3547, nx3551, 
      nx3553, nx3555, nx3559, nx3561, nx3564, nx3568, nx3572, nx3575, nx3579, 
      nx3583, nx3587, nx3589, nx3591, nx3594, nx3598, nx3602, nx3606, nx3610, 
      nx3614, nx3616, nx3618, nx3622, nx3624, nx3627, nx3632, nx3636, nx3638, 
      nx3640, nx3643, nx3648, nx3652, nx3665, nx3667, nx3669, nx3671, nx3673, 
      nx3675, nx3677, nx3679, nx3681, nx3683, nx3685, nx3687, nx3689, nx3691, 
      nx3693, nx3695, nx3697, nx3699, nx3701, nx3703, nx3705, nx3707, nx3709, 
      nx3711, nx3713, nx3715, nx3717, nx3719, nx3721, nx3723, nx3725, nx3727, 
      nx3729, nx3731, nx3733, nx3735, nx3737, nx3739, nx3741, nx3743, nx3745, 
      nx3747, nx3749, nx3751, nx3753, nx3755, nx3757, nx3759, nx3761, nx3763, 
      nx3765, nx3767, nx3769, nx3771, nx3773, nx3775, nx3777, nx3779, nx3781, 
      nx3783, nx3785, nx3787, nx3789, nx3791: std_logic ;

begin
   Product(0) <= Product_0_EXMPLR ;
   ix2791 : xor2 port map ( Y=>Product(15), A0=>nx1094, A1=>nx1260);
   ix1095 : nor02ii port map ( Y=>nx1094, A0=>nx1551, A1=>nx938);
   ix1552 : xnor2 port map ( Y=>nx1551, A0=>nx1553, A1=>nx2301);
   ix1554 : aoi32 port map ( Y=>nx1553, A0=>nx3737, A1=>nx3725, A2=>nx932, 
      B0=>nx800, B1=>nx934);
   ix933 : xnor2 port map ( Y=>nx932, A0=>nx808, A1=>nx2093);
   ix809 : oai32 port map ( Y=>nx808, A0=>nx1559, A1=>nx1561, A2=>nx1563, B0
      =>nx2005, B1=>nx2089);
   ix1560 : inv01 port map ( Y=>nx1559, A=>B(11));
   ix1562 : inv01 port map ( Y=>nx1561, A=>A(1));
   ix1564 : xnor2 port map ( Y=>nx1563, A0=>nx684, A1=>nx782);
   ix685 : oai32 port map ( Y=>nx684, A0=>nx1567, A1=>nx1569, A2=>nx1571, B0
      =>nx1851, B1=>nx1921);
   ix1568 : inv01 port map ( Y=>nx1567, A=>B(9));
   ix1570 : inv01 port map ( Y=>nx1569, A=>A(2));
   ix1572 : xnor2 port map ( Y=>nx1571, A0=>nx1573, A1=>nx1787);
   ix1574 : aoi32 port map ( Y=>nx1573, A0=>nx3761, A1=>nx3713, A2=>nx524, 
      B0=>nx464, B1=>nx526);
   ix525 : xnor2 port map ( Y=>nx524, A0=>nx472, A1=>nx1683);
   ix473 : oai32 port map ( Y=>nx472, A0=>nx1579, A1=>nx1581, A2=>nx1583, B0
      =>nx1647, B1=>nx1679);
   ix1580 : inv02 port map ( Y=>nx1579, A=>B(5));
   ix1582 : inv02 port map ( Y=>nx1581, A=>A(4));
   ix1584 : xnor2 port map ( Y=>nx1583, A0=>nx384, A1=>nx410);
   ix385 : oai32 port map ( Y=>nx384, A0=>nx1587, A1=>nx1589, A2=>nx1591, B0
      =>nx1601, B1=>nx1615);
   ix1588 : inv02 port map ( Y=>nx1587, A=>B(3));
   ix1590 : inv01 port map ( Y=>nx1589, A=>A(5));
   ix1592 : xnor2 port map ( Y=>nx1591, A0=>nx1593, A1=>nx1595);
   ix1594 : nand02 port map ( Y=>nx1593, A0=>nx3781, A1=>nx3701);
   ix1596 : xnor2 port map ( Y=>nx1595, A0=>nx1597, A1=>nx1599);
   ix1598 : nand02 port map ( Y=>nx1597, A0=>nx3785, A1=>nx3697);
   ix1600 : nand02 port map ( Y=>nx1599, A0=>nx3693, A1=>nx3789);
   ix1606 : inv01 port map ( Y=>nx1605, A=>A(7));
   ix1608 : inv01 port map ( Y=>nx1607, A=>B(0));
   ix1612 : nand02 port map ( Y=>nx1611, A0=>nx3785, A1=>nx3701);
   ix1614 : nand02 port map ( Y=>nx1613, A0=>nx3697, A1=>nx3789);
   ix1616 : xnor2 port map ( Y=>nx1615, A0=>nx1617, A1=>nx1591);
   ix1618 : nand02 port map ( Y=>nx1617, A0=>nx3777, A1=>nx3705);
   ix411 : xnor2 port map ( Y=>nx410, A0=>nx1621, A1=>nx408);
   ix1622 : nand02 port map ( Y=>nx1621, A0=>nx3773, A1=>nx3705);
   ix409 : xnor2 port map ( Y=>nx408, A0=>nx392, A1=>nx1633);
   ix393 : oai33 port map ( Y=>nx392, A0=>nx1627, A1=>nx1629, A2=>nx1595, B0
      =>nx1631, B1=>nx1605, B2=>nx1599);
   ix1628 : inv02 port map ( Y=>nx1627, A=>B(2));
   ix1630 : inv01 port map ( Y=>nx1629, A=>A(6));
   ix1632 : inv02 port map ( Y=>nx1631, A=>B(1));
   ix1634 : xnor2 port map ( Y=>nx1633, A0=>nx1635, A1=>nx1637);
   ix1636 : nand02 port map ( Y=>nx1635, A0=>nx3777, A1=>nx3701);
   ix1638 : xnor2 port map ( Y=>nx1637, A0=>nx1639, A1=>nx1641);
   ix1640 : nand02 port map ( Y=>nx1639, A0=>nx3781, A1=>nx3697);
   ix1642 : xnor2 port map ( Y=>nx1641, A0=>nx1643, A1=>nx1645);
   ix1644 : nand02 port map ( Y=>nx1643, A0=>nx3785, A1=>nx3693);
   ix1646 : nand02 port map ( Y=>nx1645, A0=>nx3689, A1=>nx3789);
   ix1648 : aoi32 port map ( Y=>nx1647, A0=>nx3773, A1=>nx3709, A2=>nx316, 
      B0=>nx292, B1=>nx318);
   ix317 : xnor2 port map ( Y=>nx316, A0=>nx300, A1=>nx1615);
   ix301 : oai33 port map ( Y=>nx300, A0=>nx1627, A1=>nx1589, A2=>nx1653, B0
      =>nx1631, B1=>nx1629, B2=>nx1613);
   ix1654 : xnor2 port map ( Y=>nx1653, A0=>nx1611, A1=>nx1613);
   ix293 : oai32 port map ( Y=>nx292, A0=>nx1587, A1=>nx1581, A2=>nx1657, B0
      =>nx1661, B1=>nx1671);
   ix1658 : xnor2 port map ( Y=>nx1657, A0=>nx1659, A1=>nx1653);
   ix1660 : nand02 port map ( Y=>nx1659, A0=>nx3781, A1=>nx3705);
   ix1668 : nand02 port map ( Y=>nx1667, A0=>nx3785, A1=>nx3705);
   ix1670 : nand02 port map ( Y=>nx1669, A0=>nx3701, A1=>nx3789);
   ix1672 : xnor2 port map ( Y=>nx1671, A0=>nx1673, A1=>nx1657);
   ix1674 : nand02 port map ( Y=>nx1673, A0=>nx3777, A1=>nx3709);
   ix319 : xnor2 port map ( Y=>nx318, A0=>nx1677, A1=>nx316);
   ix1678 : nand02 port map ( Y=>nx1677, A0=>nx3773, A1=>nx3709);
   ix1680 : xnor2 port map ( Y=>nx1679, A0=>nx1681, A1=>nx1583);
   ix1682 : nand02 port map ( Y=>nx1681, A0=>nx3769, A1=>nx3709);
   ix1684 : xnor2 port map ( Y=>nx1683, A0=>nx1685, A1=>nx1687);
   ix1686 : nand02 port map ( Y=>nx1685, A0=>nx3765, A1=>nx3709);
   ix1688 : xnor2 port map ( Y=>nx1687, A0=>nx1689, A1=>nx1691);
   ix1690 : aoi32 port map ( Y=>nx1689, A0=>nx3773, A1=>nx3705, A2=>nx408, 
      B0=>nx384, B1=>nx410);
   ix1692 : xnor2 port map ( Y=>nx1691, A0=>nx1693, A1=>nx1695);
   ix1694 : nand02 port map ( Y=>nx1693, A0=>nx3769, A1=>nx3705);
   ix1696 : xnor2 port map ( Y=>nx1695, A0=>nx488, A1=>nx514);
   ix489 : oai32 port map ( Y=>nx488, A0=>nx1587, A1=>nx1629, A2=>nx1637, B0
      =>nx1699, B1=>nx1633);
   ix1704 : inv01 port map ( Y=>nx1703, A=>A(8));
   ix515 : xnor2 port map ( Y=>nx514, A0=>nx1709, A1=>nx512);
   ix1710 : nand02 port map ( Y=>nx1709, A0=>nx3773, A1=>nx3701);
   ix513 : xnor2 port map ( Y=>nx512, A0=>nx496, A1=>nx1715);
   ix497 : oai33 port map ( Y=>nx496, A0=>nx1627, A1=>nx1605, A2=>nx1641, B0
      =>nx1631, B1=>nx1703, B2=>nx1645);
   ix1716 : xnor2 port map ( Y=>nx1715, A0=>nx1717, A1=>nx1719);
   ix1718 : nand02 port map ( Y=>nx1717, A0=>nx3777, A1=>nx3697);
   ix1720 : xnor2 port map ( Y=>nx1719, A0=>nx1721, A1=>nx1723);
   ix1722 : nand02 port map ( Y=>nx1721, A0=>nx3781, A1=>nx3693);
   ix1724 : xnor2 port map ( Y=>nx1723, A0=>nx1725, A1=>nx1727);
   ix1726 : nand02 port map ( Y=>nx1725, A0=>nx3785, A1=>nx3689);
   ix1728 : nand02 port map ( Y=>nx1727, A0=>nx3685, A1=>nx3789);
   ix465 : oai32 port map ( Y=>nx464, A0=>nx1731, A1=>nx1733, A2=>nx1735, B0
      =>nx1737, B1=>nx1779);
   ix1732 : inv02 port map ( Y=>nx1731, A=>B(6));
   ix1734 : inv01 port map ( Y=>nx1733, A=>A(3));
   ix1736 : xnor2 port map ( Y=>nx1735, A0=>nx1647, A1=>nx1679);
   ix1738 : inv01 port map ( Y=>nx1737, A=>nx368);
   ix369 : oai32 port map ( Y=>nx368, A0=>nx1579, A1=>nx1733, A2=>nx1741, B0
      =>nx1743, B1=>nx1775);
   ix1742 : xnor2 port map ( Y=>nx1741, A0=>nx292, A1=>nx318);
   ix1744 : aoi32 port map ( Y=>nx1743, A0=>nx3773, A1=>nx3713, A2=>nx236, 
      B0=>nx212, B1=>nx238);
   ix237 : xnor2 port map ( Y=>nx236, A0=>nx220, A1=>nx1671);
   ix221 : oai33 port map ( Y=>nx220, A0=>nx1627, A1=>nx1581, A2=>nx1749, B0
      =>nx1631, B1=>nx1589, B2=>nx1669);
   ix1750 : xnor2 port map ( Y=>nx1749, A0=>nx1667, A1=>nx1669);
   ix213 : oai32 port map ( Y=>nx212, A0=>nx1587, A1=>nx1733, A2=>nx1753, B0
      =>nx1757, B1=>nx1767);
   ix1754 : xnor2 port map ( Y=>nx1753, A0=>nx1755, A1=>nx1749);
   ix1756 : nand02 port map ( Y=>nx1755, A0=>nx3781, A1=>nx3709);
   ix1764 : nand02 port map ( Y=>nx1763, A0=>nx3785, A1=>nx3709);
   ix1766 : nand02 port map ( Y=>nx1765, A0=>nx3705, A1=>nx3789);
   ix1768 : xnor2 port map ( Y=>nx1767, A0=>nx1769, A1=>nx1753);
   ix1770 : nand02 port map ( Y=>nx1769, A0=>nx3777, A1=>nx3713);
   ix239 : xnor2 port map ( Y=>nx238, A0=>nx1773, A1=>nx236);
   ix1774 : nand02 port map ( Y=>nx1773, A0=>nx3773, A1=>nx3713);
   ix1776 : xnor2 port map ( Y=>nx1775, A0=>nx1777, A1=>nx1741);
   ix1778 : nand02 port map ( Y=>nx1777, A0=>nx3769, A1=>nx3713);
   ix1780 : xnor2 port map ( Y=>nx1779, A0=>nx1781, A1=>nx1735);
   ix1782 : nand02 port map ( Y=>nx1781, A0=>nx3765, A1=>nx3713);
   ix527 : xnor2 port map ( Y=>nx526, A0=>nx1785, A1=>nx524);
   ix1786 : nand02 port map ( Y=>nx1785, A0=>nx3761, A1=>nx3713);
   ix1788 : xnor2 port map ( Y=>nx1787, A0=>nx1789, A1=>nx1791);
   ix1790 : nand02 port map ( Y=>nx1789, A0=>nx3757, A1=>nx3713);
   ix1792 : xnor2 port map ( Y=>nx1791, A0=>nx580, A1=>nx642);
   ix581 : oai32 port map ( Y=>nx580, A0=>nx1731, A1=>nx1581, A2=>nx1687, B0
      =>nx1795, B1=>nx1683);
   ix1796 : inv01 port map ( Y=>nx1795, A=>nx472);
   ix643 : xnor2 port map ( Y=>nx642, A0=>nx1799, A1=>nx640);
   ix1800 : nand02 port map ( Y=>nx1799, A0=>nx3761, A1=>nx3709);
   ix641 : xnor2 port map ( Y=>nx640, A0=>nx588, A1=>nx1805);
   ix589 : oai32 port map ( Y=>nx588, A0=>nx1579, A1=>nx1589, A2=>nx1695, B0
      =>nx1689, B1=>nx1691);
   ix1806 : xnor2 port map ( Y=>nx1805, A0=>nx1807, A1=>nx1809);
   ix1808 : nand02 port map ( Y=>nx1807, A0=>nx3765, A1=>nx3705);
   ix1810 : xnor2 port map ( Y=>nx1809, A0=>nx1811, A1=>nx1813);
   ix1812 : aoi32 port map ( Y=>nx1811, A0=>nx3773, A1=>nx3701, A2=>nx512, 
      B0=>nx488, B1=>nx514);
   ix1814 : xnor2 port map ( Y=>nx1813, A0=>nx1815, A1=>nx1817);
   ix1816 : nand02 port map ( Y=>nx1815, A0=>nx3769, A1=>nx3701);
   ix1818 : xnor2 port map ( Y=>nx1817, A0=>nx604, A1=>nx630);
   ix605 : oai32 port map ( Y=>nx604, A0=>nx1587, A1=>nx1605, A2=>nx1719, B0
      =>nx1821, B1=>nx1715);
   ix1826 : inv01 port map ( Y=>nx1825, A=>A(9));
   ix631 : xnor2 port map ( Y=>nx630, A0=>nx1831, A1=>nx628);
   ix1832 : nand02 port map ( Y=>nx1831, A0=>nx3773, A1=>nx3697);
   ix629 : xnor2 port map ( Y=>nx628, A0=>nx612, A1=>nx1837);
   ix613 : oai33 port map ( Y=>nx612, A0=>nx1627, A1=>nx1703, A2=>nx1723, B0
      =>nx1631, B1=>nx1825, B2=>nx1727);
   ix1838 : xnor2 port map ( Y=>nx1837, A0=>nx1839, A1=>nx1841);
   ix1840 : nand02 port map ( Y=>nx1839, A0=>nx3777, A1=>nx3693);
   ix1842 : xnor2 port map ( Y=>nx1841, A0=>nx1843, A1=>nx1845);
   ix1844 : nand02 port map ( Y=>nx1843, A0=>nx3781, A1=>nx3689);
   ix1846 : xnor2 port map ( Y=>nx1845, A0=>nx1847, A1=>nx1849);
   ix1848 : nand02 port map ( Y=>nx1847, A0=>nx3785, A1=>nx3685);
   ix1850 : nand02 port map ( Y=>nx1849, A0=>nx3681, A1=>nx3789);
   ix1852 : inv01 port map ( Y=>nx1851, A=>nx564);
   ix565 : oai32 port map ( Y=>nx564, A0=>nx1855, A1=>nx1569, A2=>nx1857, B0
      =>nx1859, B1=>nx1917);
   ix1856 : inv01 port map ( Y=>nx1855, A=>B(8));
   ix1858 : xnor2 port map ( Y=>nx1857, A0=>nx464, A1=>nx526);
   ix1860 : aoi32 port map ( Y=>nx1859, A0=>nx3761, A1=>nx3717, A2=>nx420, 
      B0=>nx360, B1=>nx422);
   ix421 : xnor2 port map ( Y=>nx420, A0=>nx368, A1=>nx1779);
   ix361 : oai32 port map ( Y=>nx360, A0=>nx1731, A1=>nx1569, A2=>nx1865, B0
      =>nx1867, B1=>nx1909);
   ix1866 : xnor2 port map ( Y=>nx1865, A0=>nx1743, A1=>nx1775);
   ix1868 : inv01 port map ( Y=>nx1867, A=>nx276);
   ix277 : oai32 port map ( Y=>nx276, A0=>nx1579, A1=>nx1569, A2=>nx1871, B0
      =>nx1873, B1=>nx1905);
   ix1872 : xnor2 port map ( Y=>nx1871, A0=>nx212, A1=>nx238);
   ix1874 : aoi32 port map ( Y=>nx1873, A0=>nx3773, A1=>nx3717, A2=>nx168, 
      B0=>nx144, B1=>nx170);
   ix169 : xnor2 port map ( Y=>nx168, A0=>nx152, A1=>nx1767);
   ix153 : oai33 port map ( Y=>nx152, A0=>nx1627, A1=>nx1733, A2=>nx1879, B0
      =>nx1631, B1=>nx1581, B2=>nx1765);
   ix1880 : xnor2 port map ( Y=>nx1879, A0=>nx1763, A1=>nx1765);
   ix145 : oai32 port map ( Y=>nx144, A0=>nx1587, A1=>nx1569, A2=>nx1883, B0
      =>nx1887, B1=>nx1897);
   ix1884 : xnor2 port map ( Y=>nx1883, A0=>nx1885, A1=>nx1879);
   ix1886 : nand02 port map ( Y=>nx1885, A0=>nx3781, A1=>nx3713);
   ix1894 : nand02 port map ( Y=>nx1893, A0=>nx3785, A1=>nx3713);
   ix1896 : nand02 port map ( Y=>nx1895, A0=>nx3709, A1=>nx3789);
   ix1898 : xnor2 port map ( Y=>nx1897, A0=>nx1899, A1=>nx1883);
   ix1900 : nand02 port map ( Y=>nx1899, A0=>nx3777, A1=>nx3717);
   ix171 : xnor2 port map ( Y=>nx170, A0=>nx1903, A1=>nx168);
   ix1904 : nand02 port map ( Y=>nx1903, A0=>nx3773, A1=>nx3717);
   ix1906 : xnor2 port map ( Y=>nx1905, A0=>nx1907, A1=>nx1871);
   ix1908 : nand02 port map ( Y=>nx1907, A0=>nx3769, A1=>nx3717);
   ix1910 : xnor2 port map ( Y=>nx1909, A0=>nx1911, A1=>nx1865);
   ix1912 : nand02 port map ( Y=>nx1911, A0=>nx3765, A1=>nx3717);
   ix423 : xnor2 port map ( Y=>nx422, A0=>nx1915, A1=>nx420);
   ix1916 : nand02 port map ( Y=>nx1915, A0=>nx3761, A1=>nx3717);
   ix1918 : xnor2 port map ( Y=>nx1917, A0=>nx1919, A1=>nx1857);
   ix1920 : nand02 port map ( Y=>nx1919, A0=>nx3757, A1=>nx3717);
   ix1922 : xnor2 port map ( Y=>nx1921, A0=>nx1923, A1=>nx1571);
   ix1924 : nand02 port map ( Y=>nx1923, A0=>nx3753, A1=>nx3717);
   ix783 : xnor2 port map ( Y=>nx782, A0=>nx1927, A1=>nx780);
   ix1928 : nand02 port map ( Y=>nx1927, A0=>nx3749, A1=>nx3717);
   ix781 : xnor2 port map ( Y=>nx780, A0=>nx692, A1=>nx1933);
   ix693 : oai32 port map ( Y=>nx692, A0=>nx1855, A1=>nx1733, A2=>nx1791, B0
      =>nx1573, B1=>nx1787);
   ix1934 : xnor2 port map ( Y=>nx1933, A0=>nx1935, A1=>nx1937);
   ix1936 : nand02 port map ( Y=>nx1935, A0=>nx3753, A1=>nx3713);
   ix1938 : xnor2 port map ( Y=>nx1937, A0=>nx1939, A1=>nx1941);
   ix1940 : aoi32 port map ( Y=>nx1939, A0=>nx3761, A1=>nx3709, A2=>nx640, 
      B0=>nx580, B1=>nx642);
   ix1942 : xnor2 port map ( Y=>nx1941, A0=>nx1943, A1=>nx1945);
   ix1944 : nand02 port map ( Y=>nx1943, A0=>nx3757, A1=>nx3709);
   ix1946 : xnor2 port map ( Y=>nx1945, A0=>nx708, A1=>nx770);
   ix709 : oai32 port map ( Y=>nx708, A0=>nx1731, A1=>nx1589, A2=>nx1809, B0
      =>nx1949, B1=>nx1805);
   ix1950 : inv01 port map ( Y=>nx1949, A=>nx588);
   ix771 : xnor2 port map ( Y=>nx770, A0=>nx1953, A1=>nx768);
   ix1954 : nand02 port map ( Y=>nx1953, A0=>nx3761, A1=>nx3705);
   ix769 : xnor2 port map ( Y=>nx768, A0=>nx716, A1=>nx1959);
   ix717 : oai32 port map ( Y=>nx716, A0=>nx1579, A1=>nx1629, A2=>nx1817, B0
      =>nx1811, B1=>nx1813);
   ix1960 : xnor2 port map ( Y=>nx1959, A0=>nx1961, A1=>nx1963);
   ix1962 : nand02 port map ( Y=>nx1961, A0=>nx3765, A1=>nx3701);
   ix1964 : xnor2 port map ( Y=>nx1963, A0=>nx1965, A1=>nx1967);
   ix1966 : aoi32 port map ( Y=>nx1965, A0=>nx3773, A1=>nx3697, A2=>nx628, 
      B0=>nx604, B1=>nx630);
   ix1968 : xnor2 port map ( Y=>nx1967, A0=>nx1969, A1=>nx1971);
   ix1970 : nand02 port map ( Y=>nx1969, A0=>nx3769, A1=>nx3697);
   ix1972 : xnor2 port map ( Y=>nx1971, A0=>nx732, A1=>nx758);
   ix733 : oai32 port map ( Y=>nx732, A0=>nx1587, A1=>nx1703, A2=>nx1841, B0
      =>nx1975, B1=>nx1837);
   ix1980 : inv01 port map ( Y=>nx1979, A=>A(10));
   ix759 : xnor2 port map ( Y=>nx758, A0=>nx1985, A1=>nx756);
   ix1986 : nand02 port map ( Y=>nx1985, A0=>nx3773, A1=>nx3693);
   ix757 : xnor2 port map ( Y=>nx756, A0=>nx740, A1=>nx1991);
   ix741 : oai33 port map ( Y=>nx740, A0=>nx1627, A1=>nx1825, A2=>nx1845, B0
      =>nx1631, B1=>nx1979, B2=>nx1849);
   ix1992 : xnor2 port map ( Y=>nx1991, A0=>nx1993, A1=>nx1995);
   ix1994 : nand02 port map ( Y=>nx1993, A0=>nx3777, A1=>nx3689);
   ix1996 : xnor2 port map ( Y=>nx1995, A0=>nx1997, A1=>nx1999);
   ix1998 : nand02 port map ( Y=>nx1997, A0=>nx3781, A1=>nx3685);
   ix2000 : xnor2 port map ( Y=>nx1999, A0=>nx2001, A1=>nx2003);
   ix2002 : nand02 port map ( Y=>nx2001, A0=>nx3785, A1=>nx3681);
   ix2004 : nand02 port map ( Y=>nx2003, A0=>nx3677, A1=>nx3789);
   ix2006 : aoi32 port map ( Y=>nx2005, A0=>nx3749, A1=>nx3721, A2=>nx652, 
      B0=>nx556, B1=>nx654);
   ix653 : xnor2 port map ( Y=>nx652, A0=>nx564, A1=>nx1921);
   ix557 : oai32 port map ( Y=>nx556, A0=>nx1567, A1=>nx1561, A2=>nx2011, B0
      =>nx2013, B1=>nx2081);
   ix2012 : xnor2 port map ( Y=>nx2011, A0=>nx1859, A1=>nx1917);
   ix2014 : inv01 port map ( Y=>nx2013, A=>nx448);
   ix449 : oai32 port map ( Y=>nx448, A0=>nx1855, A1=>nx1561, A2=>nx2017, B0
      =>nx2019, B1=>nx2077);
   ix2018 : xnor2 port map ( Y=>nx2017, A0=>nx360, A1=>nx422);
   ix2020 : aoi32 port map ( Y=>nx2019, A0=>nx3761, A1=>nx3721, A2=>nx328, 
      B0=>nx268, B1=>nx330);
   ix329 : xnor2 port map ( Y=>nx328, A0=>nx276, A1=>nx1909);
   ix269 : oai32 port map ( Y=>nx268, A0=>nx1731, A1=>nx1561, A2=>nx2025, B0
      =>nx2027, B1=>nx2069);
   ix2026 : xnor2 port map ( Y=>nx2025, A0=>nx1873, A1=>nx1905);
   ix2028 : inv01 port map ( Y=>nx2027, A=>nx196);
   ix197 : oai32 port map ( Y=>nx196, A0=>nx1579, A1=>nx1561, A2=>nx2031, B0
      =>nx2033, B1=>nx2065);
   ix2032 : xnor2 port map ( Y=>nx2031, A0=>nx144, A1=>nx170);
   ix2034 : aoi32 port map ( Y=>nx2033, A0=>nx3773, A1=>nx3721, A2=>nx112, 
      B0=>nx88, B1=>nx114);
   ix113 : xnor2 port map ( Y=>nx112, A0=>nx96, A1=>nx1897);
   ix97 : oai33 port map ( Y=>nx96, A0=>nx1627, A1=>nx1569, A2=>nx2039, B0=>
      nx1631, B1=>nx1733, B2=>nx1895);
   ix2040 : xnor2 port map ( Y=>nx2039, A0=>nx1893, A1=>nx1895);
   ix89 : oai32 port map ( Y=>nx88, A0=>nx1587, A1=>nx1561, A2=>nx2043, B0=>
      nx2047, B1=>nx2057);
   ix2044 : xnor2 port map ( Y=>nx2043, A0=>nx2045, A1=>nx2039);
   ix2046 : nand02 port map ( Y=>nx2045, A0=>nx3781, A1=>nx3717);
   ix2054 : nand02 port map ( Y=>nx2053, A0=>nx3785, A1=>nx3717);
   ix2056 : nand02 port map ( Y=>nx2055, A0=>nx3713, A1=>nx3789);
   ix2058 : xnor2 port map ( Y=>nx2057, A0=>nx2059, A1=>nx2043);
   ix2060 : nand02 port map ( Y=>nx2059, A0=>nx3777, A1=>nx3721);
   ix115 : xnor2 port map ( Y=>nx114, A0=>nx2063, A1=>nx112);
   ix2064 : nand02 port map ( Y=>nx2063, A0=>nx3773, A1=>nx3721);
   ix2066 : xnor2 port map ( Y=>nx2065, A0=>nx2067, A1=>nx2031);
   ix2068 : nand02 port map ( Y=>nx2067, A0=>nx3769, A1=>nx3721);
   ix2070 : xnor2 port map ( Y=>nx2069, A0=>nx2071, A1=>nx2025);
   ix2072 : nand02 port map ( Y=>nx2071, A0=>nx3765, A1=>nx3721);
   ix331 : xnor2 port map ( Y=>nx330, A0=>nx2075, A1=>nx328);
   ix2076 : nand02 port map ( Y=>nx2075, A0=>nx3761, A1=>nx3721);
   ix2078 : xnor2 port map ( Y=>nx2077, A0=>nx2079, A1=>nx2017);
   ix2080 : nand02 port map ( Y=>nx2079, A0=>nx3757, A1=>nx3721);
   ix2082 : xnor2 port map ( Y=>nx2081, A0=>nx2083, A1=>nx2011);
   ix2084 : nand02 port map ( Y=>nx2083, A0=>nx3753, A1=>nx3721);
   ix655 : xnor2 port map ( Y=>nx654, A0=>nx2087, A1=>nx652);
   ix2088 : nand02 port map ( Y=>nx2087, A0=>nx3749, A1=>nx3721);
   ix2090 : xnor2 port map ( Y=>nx2089, A0=>nx2091, A1=>nx1563);
   ix2092 : nand02 port map ( Y=>nx2091, A0=>nx3745, A1=>nx3721);
   ix2094 : xnor2 port map ( Y=>nx2093, A0=>nx2095, A1=>nx2097);
   ix2096 : nand02 port map ( Y=>nx2095, A0=>nx3741, A1=>nx3721);
   ix2098 : xnor2 port map ( Y=>nx2097, A0=>nx2099, A1=>nx2101);
   ix2100 : aoi32 port map ( Y=>nx2099, A0=>nx3749, A1=>nx3717, A2=>nx780, 
      B0=>nx684, B1=>nx782);
   ix2102 : xnor2 port map ( Y=>nx2101, A0=>nx2103, A1=>nx2105);
   ix2104 : nand02 port map ( Y=>nx2103, A0=>nx3745, A1=>nx3717);
   ix2106 : xnor2 port map ( Y=>nx2105, A0=>nx824, A1=>nx922);
   ix825 : oai32 port map ( Y=>nx824, A0=>nx1567, A1=>nx1733, A2=>nx1937, B0
      =>nx2109, B1=>nx1933);
   ix2110 : inv01 port map ( Y=>nx2109, A=>nx692);
   ix923 : xnor2 port map ( Y=>nx922, A0=>nx2113, A1=>nx920);
   ix2114 : nand02 port map ( Y=>nx2113, A0=>nx3749, A1=>nx3713);
   ix921 : xnor2 port map ( Y=>nx920, A0=>nx832, A1=>nx2119);
   ix833 : oai32 port map ( Y=>nx832, A0=>nx1855, A1=>nx1581, A2=>nx1945, B0
      =>nx1939, B1=>nx1941);
   ix2120 : xnor2 port map ( Y=>nx2119, A0=>nx2121, A1=>nx2123);
   ix2122 : nand02 port map ( Y=>nx2121, A0=>nx3753, A1=>nx3709);
   ix2124 : xnor2 port map ( Y=>nx2123, A0=>nx2125, A1=>nx2127);
   ix2126 : aoi32 port map ( Y=>nx2125, A0=>nx3761, A1=>nx3705, A2=>nx768, 
      B0=>nx708, B1=>nx770);
   ix2128 : xnor2 port map ( Y=>nx2127, A0=>nx2129, A1=>nx2131);
   ix2130 : nand02 port map ( Y=>nx2129, A0=>nx3757, A1=>nx3705);
   ix2132 : xnor2 port map ( Y=>nx2131, A0=>nx848, A1=>nx910);
   ix849 : oai32 port map ( Y=>nx848, A0=>nx1731, A1=>nx1629, A2=>nx1963, B0
      =>nx2135, B1=>nx1959);
   ix2136 : inv01 port map ( Y=>nx2135, A=>nx716);
   ix911 : xnor2 port map ( Y=>nx910, A0=>nx2139, A1=>nx908);
   ix2140 : nand02 port map ( Y=>nx2139, A0=>nx3761, A1=>nx3701);
   ix909 : xnor2 port map ( Y=>nx908, A0=>nx856, A1=>nx2145);
   ix857 : oai32 port map ( Y=>nx856, A0=>nx1579, A1=>nx1605, A2=>nx1971, B0
      =>nx1965, B1=>nx1967);
   ix2146 : xnor2 port map ( Y=>nx2145, A0=>nx2147, A1=>nx2149);
   ix2148 : nand02 port map ( Y=>nx2147, A0=>nx3765, A1=>nx3697);
   ix2150 : xnor2 port map ( Y=>nx2149, A0=>nx2151, A1=>nx2153);
   ix2152 : aoi32 port map ( Y=>nx2151, A0=>nx3775, A1=>nx3693, A2=>nx756, 
      B0=>nx732, B1=>nx758);
   ix2154 : xnor2 port map ( Y=>nx2153, A0=>nx2155, A1=>nx2157);
   ix2156 : nand02 port map ( Y=>nx2155, A0=>nx3769, A1=>nx3693);
   ix2158 : xnor2 port map ( Y=>nx2157, A0=>nx872, A1=>nx898);
   ix873 : oai32 port map ( Y=>nx872, A0=>nx1587, A1=>nx1825, A2=>nx1995, B0
      =>nx2161, B1=>nx1991);
   ix2166 : inv01 port map ( Y=>nx2165, A=>A(11));
   ix899 : xnor2 port map ( Y=>nx898, A0=>nx2171, A1=>nx896);
   ix2172 : nand02 port map ( Y=>nx2171, A0=>nx3775, A1=>nx3689);
   ix897 : xnor2 port map ( Y=>nx896, A0=>nx880, A1=>nx2177);
   ix881 : oai33 port map ( Y=>nx880, A0=>nx1627, A1=>nx1979, A2=>nx1999, B0
      =>nx1631, B1=>nx2165, B2=>nx2003);
   ix2178 : xnor2 port map ( Y=>nx2177, A0=>nx2179, A1=>nx2181);
   ix2180 : nand02 port map ( Y=>nx2179, A0=>nx3777, A1=>nx3685);
   ix2182 : xnor2 port map ( Y=>nx2181, A0=>nx2183, A1=>nx2185);
   ix2184 : nand02 port map ( Y=>nx2183, A0=>nx3781, A1=>nx3681);
   ix2186 : xnor2 port map ( Y=>nx2185, A0=>nx2187, A1=>nx2189);
   ix2188 : nand02 port map ( Y=>nx2187, A0=>nx3785, A1=>nx3677);
   ix2190 : nand02 port map ( Y=>nx2189, A0=>nx3673, A1=>nx3789);
   ix801 : oai32 port map ( Y=>nx800, A0=>nx2193, A1=>nx2195, A2=>nx2197, B0
      =>nx2199, B1=>nx2293);
   ix2194 : inv01 port map ( Y=>nx2193, A=>B(12));
   ix2196 : inv01 port map ( Y=>nx2195, A=>A(0));
   ix2198 : xnor2 port map ( Y=>nx2197, A0=>nx2005, A1=>nx2089);
   ix2200 : inv01 port map ( Y=>nx2199, A=>nx668);
   ix669 : oai32 port map ( Y=>nx668, A0=>nx1559, A1=>nx2195, A2=>nx2203, B0
      =>nx2205, B1=>nx2289);
   ix2204 : xnor2 port map ( Y=>nx2203, A0=>nx556, A1=>nx654);
   ix2206 : aoi32 port map ( Y=>nx2205, A0=>nx3749, A1=>nx3725, A2=>nx536, 
      B0=>nx440, B1=>nx538);
   ix537 : xnor2 port map ( Y=>nx536, A0=>nx448, A1=>nx2081);
   ix441 : oai32 port map ( Y=>nx440, A0=>nx1567, A1=>nx2195, A2=>nx2211, B0
      =>nx2213, B1=>nx2281);
   ix2212 : xnor2 port map ( Y=>nx2211, A0=>nx2019, A1=>nx2077);
   ix2214 : inv01 port map ( Y=>nx2213, A=>nx344);
   ix345 : oai32 port map ( Y=>nx344, A0=>nx1855, A1=>nx2195, A2=>nx2217, B0
      =>nx2219, B1=>nx2277);
   ix2218 : xnor2 port map ( Y=>nx2217, A0=>nx268, A1=>nx330);
   ix2220 : aoi32 port map ( Y=>nx2219, A0=>nx3761, A1=>nx3725, A2=>nx248, 
      B0=>nx188, B1=>nx250);
   ix249 : xnor2 port map ( Y=>nx248, A0=>nx196, A1=>nx2069);
   ix189 : oai32 port map ( Y=>nx188, A0=>nx1731, A1=>nx2195, A2=>nx2225, B0
      =>nx2227, B1=>nx2269);
   ix2226 : xnor2 port map ( Y=>nx2225, A0=>nx2033, A1=>nx2065);
   ix2228 : inv01 port map ( Y=>nx2227, A=>nx128);
   ix129 : oai32 port map ( Y=>nx128, A0=>nx1579, A1=>nx2195, A2=>nx2231, B0
      =>nx2233, B1=>nx2265);
   ix2232 : xnor2 port map ( Y=>nx2231, A0=>nx88, A1=>nx114);
   ix2234 : aoi32 port map ( Y=>nx2233, A0=>nx3775, A1=>nx3725, A2=>nx68, B0
      =>nx44, B1=>nx70);
   ix69 : xnor2 port map ( Y=>nx68, A0=>nx52, A1=>nx2057);
   ix53 : oai33 port map ( Y=>nx52, A0=>nx1627, A1=>nx1561, A2=>nx2239, B0=>
      nx1631, B1=>nx1569, B2=>nx2055);
   ix2240 : xnor2 port map ( Y=>nx2239, A0=>nx2053, A1=>nx2055);
   ix45 : oai32 port map ( Y=>nx44, A0=>nx1587, A1=>nx2195, A2=>nx2243, B0=>
      nx2247, B1=>nx2257);
   ix2244 : xnor2 port map ( Y=>nx2243, A0=>nx2245, A1=>nx2239);
   ix2246 : nand02 port map ( Y=>nx2245, A0=>nx3781, A1=>nx3721);
   ix2254 : nand02 port map ( Y=>nx2253, A0=>nx3785, A1=>nx3721);
   ix2256 : nand02 port map ( Y=>nx2255, A0=>nx3717, A1=>nx3789);
   ix2258 : xnor2 port map ( Y=>nx2257, A0=>nx2259, A1=>nx2243);
   ix2260 : nand02 port map ( Y=>nx2259, A0=>nx3777, A1=>nx3725);
   ix71 : xnor2 port map ( Y=>nx70, A0=>nx2263, A1=>nx68);
   ix2264 : nand02 port map ( Y=>nx2263, A0=>nx3775, A1=>nx3725);
   ix2266 : xnor2 port map ( Y=>nx2265, A0=>nx2267, A1=>nx2231);
   ix2268 : nand02 port map ( Y=>nx2267, A0=>nx3769, A1=>nx3725);
   ix2270 : xnor2 port map ( Y=>nx2269, A0=>nx2271, A1=>nx2225);
   ix2272 : nand02 port map ( Y=>nx2271, A0=>nx3765, A1=>nx3725);
   ix251 : xnor2 port map ( Y=>nx250, A0=>nx2275, A1=>nx248);
   ix2276 : nand02 port map ( Y=>nx2275, A0=>nx3761, A1=>nx3725);
   ix2278 : xnor2 port map ( Y=>nx2277, A0=>nx2279, A1=>nx2217);
   ix2280 : nand02 port map ( Y=>nx2279, A0=>nx3757, A1=>nx3725);
   ix2282 : xnor2 port map ( Y=>nx2281, A0=>nx2283, A1=>nx2211);
   ix2284 : nand02 port map ( Y=>nx2283, A0=>nx3753, A1=>nx3725);
   ix539 : xnor2 port map ( Y=>nx538, A0=>nx2287, A1=>nx536);
   ix2288 : nand02 port map ( Y=>nx2287, A0=>nx3749, A1=>nx3725);
   ix2290 : xnor2 port map ( Y=>nx2289, A0=>nx2291, A1=>nx2203);
   ix2292 : nand02 port map ( Y=>nx2291, A0=>nx3745, A1=>nx3725);
   ix2294 : xnor2 port map ( Y=>nx2293, A0=>nx2295, A1=>nx2197);
   ix2296 : nand02 port map ( Y=>nx2295, A0=>nx3741, A1=>nx3725);
   ix935 : xnor2 port map ( Y=>nx934, A0=>nx2299, A1=>nx932);
   ix2300 : nand02 port map ( Y=>nx2299, A0=>nx3737, A1=>nx3725);
   ix2302 : xnor2 port map ( Y=>nx2301, A0=>nx2303, A1=>nx2305);
   ix2304 : nand02 port map ( Y=>nx2303, A0=>nx3733, A1=>nx3727);
   ix2306 : xnor2 port map ( Y=>nx2305, A0=>nx952, A1=>nx1086);
   ix953 : oai32 port map ( Y=>nx952, A0=>nx2193, A1=>nx1561, A2=>nx2097, B0
      =>nx2309, B1=>nx2093);
   ix2310 : inv01 port map ( Y=>nx2309, A=>nx808);
   ix1087 : xnor2 port map ( Y=>nx1086, A0=>nx2313, A1=>nx1084);
   ix2314 : nand02 port map ( Y=>nx2313, A0=>nx3737, A1=>nx3723);
   ix1085 : xnor2 port map ( Y=>nx1084, A0=>nx960, A1=>nx2319);
   ix961 : oai32 port map ( Y=>nx960, A0=>nx1559, A1=>nx1569, A2=>nx2105, B0
      =>nx2099, B1=>nx2101);
   ix2320 : xnor2 port map ( Y=>nx2319, A0=>nx2321, A1=>nx2323);
   ix2322 : nand02 port map ( Y=>nx2321, A0=>nx3741, A1=>nx3719);
   ix2324 : xnor2 port map ( Y=>nx2323, A0=>nx2325, A1=>nx2327);
   ix2326 : aoi32 port map ( Y=>nx2325, A0=>nx3749, A1=>nx3713, A2=>nx920, 
      B0=>nx824, B1=>nx922);
   ix2328 : xnor2 port map ( Y=>nx2327, A0=>nx2329, A1=>nx2331);
   ix2330 : nand02 port map ( Y=>nx2329, A0=>nx3745, A1=>nx3713);
   ix2332 : xnor2 port map ( Y=>nx2331, A0=>nx976, A1=>nx1074);
   ix977 : oai32 port map ( Y=>nx976, A0=>nx1567, A1=>nx1581, A2=>nx2123, B0
      =>nx2335, B1=>nx2119);
   ix2336 : inv01 port map ( Y=>nx2335, A=>nx832);
   ix1075 : xnor2 port map ( Y=>nx1074, A0=>nx2339, A1=>nx1072);
   ix2340 : nand02 port map ( Y=>nx2339, A0=>nx3749, A1=>nx3709);
   ix1073 : xnor2 port map ( Y=>nx1072, A0=>nx984, A1=>nx2345);
   ix985 : oai32 port map ( Y=>nx984, A0=>nx1855, A1=>nx1589, A2=>nx2131, B0
      =>nx2125, B1=>nx2127);
   ix2346 : xnor2 port map ( Y=>nx2345, A0=>nx2347, A1=>nx2349);
   ix2348 : nand02 port map ( Y=>nx2347, A0=>nx3753, A1=>nx3705);
   ix2350 : xnor2 port map ( Y=>nx2349, A0=>nx2351, A1=>nx2353);
   ix2352 : aoi32 port map ( Y=>nx2351, A0=>nx3761, A1=>nx3701, A2=>nx908, 
      B0=>nx848, B1=>nx910);
   ix2354 : xnor2 port map ( Y=>nx2353, A0=>nx2355, A1=>nx2357);
   ix2356 : nand02 port map ( Y=>nx2355, A0=>nx3757, A1=>nx3701);
   ix2358 : xnor2 port map ( Y=>nx2357, A0=>nx1000, A1=>nx1062);
   ix1001 : oai32 port map ( Y=>nx1000, A0=>nx1731, A1=>nx1605, A2=>nx2149, 
      B0=>nx2361, B1=>nx2145);
   ix2362 : inv01 port map ( Y=>nx2361, A=>nx856);
   ix1063 : xnor2 port map ( Y=>nx1062, A0=>nx2365, A1=>nx1060);
   ix2366 : nand02 port map ( Y=>nx2365, A0=>nx3761, A1=>nx3697);
   ix1061 : xnor2 port map ( Y=>nx1060, A0=>nx1008, A1=>nx2371);
   ix1009 : oai32 port map ( Y=>nx1008, A0=>nx1579, A1=>nx1703, A2=>nx2157, 
      B0=>nx2151, B1=>nx2153);
   ix2372 : xnor2 port map ( Y=>nx2371, A0=>nx2373, A1=>nx2375);
   ix2374 : nand02 port map ( Y=>nx2373, A0=>nx3765, A1=>nx3693);
   ix2376 : xnor2 port map ( Y=>nx2375, A0=>nx2377, A1=>nx2379);
   ix2378 : aoi32 port map ( Y=>nx2377, A0=>nx3775, A1=>nx3689, A2=>nx896, 
      B0=>nx872, B1=>nx898);
   ix2380 : xnor2 port map ( Y=>nx2379, A0=>nx2381, A1=>nx2383);
   ix2382 : nand02 port map ( Y=>nx2381, A0=>nx3769, A1=>nx3689);
   ix2384 : xnor2 port map ( Y=>nx2383, A0=>nx1024, A1=>nx1050);
   ix1025 : oai32 port map ( Y=>nx1024, A0=>nx1587, A1=>nx1979, A2=>nx2181, 
      B0=>nx2387, B1=>nx2177);
   ix2392 : inv01 port map ( Y=>nx2391, A=>A(12));
   ix1051 : xnor2 port map ( Y=>nx1050, A0=>nx2397, A1=>nx1048);
   ix2398 : nand02 port map ( Y=>nx2397, A0=>nx3775, A1=>nx3685);
   ix1049 : xnor2 port map ( Y=>nx1048, A0=>nx1032, A1=>nx2403);
   ix1033 : oai33 port map ( Y=>nx1032, A0=>nx1627, A1=>nx2165, A2=>nx2185, 
      B0=>nx1631, B1=>nx2391, B2=>nx2189);
   ix2404 : xnor2 port map ( Y=>nx2403, A0=>nx2405, A1=>nx2407);
   ix2406 : nand02 port map ( Y=>nx2405, A0=>nx3777, A1=>nx3681);
   ix2408 : xnor2 port map ( Y=>nx2407, A0=>nx2409, A1=>nx2411);
   ix2410 : nand02 port map ( Y=>nx2409, A0=>nx3781, A1=>nx3677);
   ix2412 : xnor2 port map ( Y=>nx2411, A0=>nx2413, A1=>nx2415);
   ix2414 : nand02 port map ( Y=>nx2413, A0=>nx3785, A1=>nx3673);
   ix2416 : nand02 port map ( Y=>nx2415, A0=>nx3669, A1=>nx3789);
   ix939 : nor02 port map ( Y=>nx938, A0=>nx2419, A1=>nx2473);
   ix2420 : nand02 port map ( Y=>nx2419, A0=>nx662, A1=>nx792);
   ix663 : nor02ii port map ( Y=>nx662, A0=>nx2423, A1=>nx542);
   ix2424 : xnor2 port map ( Y=>nx2423, A0=>nx2205, A1=>nx2289);
   ix543 : nor02 port map ( Y=>nx542, A0=>nx2427, A1=>nx2469);
   ix2428 : nand02 port map ( Y=>nx2427, A0=>nx338, A1=>nx432);
   ix339 : nor02ii port map ( Y=>nx338, A0=>nx2431, A1=>nx254);
   ix2432 : xnor2 port map ( Y=>nx2431, A0=>nx2219, A1=>nx2277);
   ix255 : nor02 port map ( Y=>nx254, A0=>nx2435, A1=>nx2465);
   ix2436 : nand02 port map ( Y=>nx2435, A0=>nx122, A1=>nx180);
   ix123 : nor02ii port map ( Y=>nx122, A0=>nx2439, A1=>nx74);
   ix2440 : xnor2 port map ( Y=>nx2439, A0=>nx2233, A1=>nx2265);
   ix75 : nor02 port map ( Y=>nx74, A0=>nx2443, A1=>nx2461);
   ix2444 : nand02 port map ( Y=>nx2443, A0=>nx14, A1=>nx36);
   ix15 : nor02 port map ( Y=>nx14, A0=>nx2447, A1=>nx2451);
   ix2448 : nand03 port map ( Y=>nx2447, A0=>nx3785, A1=>nx3723, A2=>
      Product_0_EXMPLR);
   ix2452 : xnor2 port map ( Y=>nx2451, A0=>nx2453, A1=>nx2455);
   ix2454 : nand02 port map ( Y=>nx2453, A0=>nx3781, A1=>nx3727);
   ix2456 : xnor2 port map ( Y=>nx2455, A0=>nx2253, A1=>nx2255);
   ix37 : xnor2 port map ( Y=>nx36, A0=>nx20, A1=>nx2257);
   ix21 : oai33 port map ( Y=>nx20, A0=>nx1627, A1=>nx2195, A2=>nx2455, B0=>
      nx2253, B1=>nx1569, B2=>nx1607);
   ix2462 : xnor2 port map ( Y=>nx2461, A0=>nx44, A1=>nx70);
   ix181 : xnor2 port map ( Y=>nx180, A0=>nx128, A1=>nx2269);
   ix2466 : xnor2 port map ( Y=>nx2465, A0=>nx188, A1=>nx250);
   ix433 : xnor2 port map ( Y=>nx432, A0=>nx344, A1=>nx2281);
   ix2470 : xnor2 port map ( Y=>nx2469, A0=>nx440, A1=>nx538);
   ix793 : xnor2 port map ( Y=>nx792, A0=>nx668, A1=>nx2293);
   ix2474 : xnor2 port map ( Y=>nx2473, A0=>nx800, A1=>nx934);
   ix1261 : xnor2 port map ( Y=>nx1260, A0=>nx1100, A1=>nx2481);
   ix1101 : oai32 port map ( Y=>nx1100, A0=>nx2479, A1=>nx2195, A2=>nx2305, 
      B0=>nx1553, B1=>nx2301);
   ix2480 : inv01 port map ( Y=>nx2479, A=>B(14));
   ix2482 : xnor2 port map ( Y=>nx2481, A0=>nx2483, A1=>nx2485);
   ix2484 : nand02 port map ( Y=>nx2483, A0=>nx3729, A1=>nx3727);
   ix2486 : xnor2 port map ( Y=>nx2485, A0=>nx2487, A1=>nx2489);
   ix2488 : aoi32 port map ( Y=>nx2487, A0=>nx3737, A1=>nx3723, A2=>nx1084, 
      B0=>nx952, B1=>nx1086);
   ix2490 : xnor2 port map ( Y=>nx2489, A0=>nx2491, A1=>nx2493);
   ix2492 : nand02 port map ( Y=>nx2491, A0=>nx3733, A1=>nx3723);
   ix2494 : xnor2 port map ( Y=>nx2493, A0=>nx1116, A1=>nx1250);
   ix1117 : oai32 port map ( Y=>nx1116, A0=>nx2193, A1=>nx1569, A2=>nx2323, 
      B0=>nx2497, B1=>nx2319);
   ix2498 : inv01 port map ( Y=>nx2497, A=>nx960);
   ix1251 : xnor2 port map ( Y=>nx1250, A0=>nx2501, A1=>nx1248);
   ix2502 : nand02 port map ( Y=>nx2501, A0=>nx3737, A1=>nx3719);
   ix1249 : xnor2 port map ( Y=>nx1248, A0=>nx1124, A1=>nx2507);
   ix1125 : oai32 port map ( Y=>nx1124, A0=>nx1559, A1=>nx1733, A2=>nx2331, 
      B0=>nx2325, B1=>nx2327);
   ix2508 : xnor2 port map ( Y=>nx2507, A0=>nx2509, A1=>nx2511);
   ix2510 : nand02 port map ( Y=>nx2509, A0=>nx3741, A1=>nx3715);
   ix2512 : xnor2 port map ( Y=>nx2511, A0=>nx2513, A1=>nx2515);
   ix2514 : aoi32 port map ( Y=>nx2513, A0=>nx3749, A1=>nx3709, A2=>nx1072, 
      B0=>nx976, B1=>nx1074);
   ix2516 : xnor2 port map ( Y=>nx2515, A0=>nx2517, A1=>nx2519);
   ix2518 : nand02 port map ( Y=>nx2517, A0=>nx3745, A1=>nx3709);
   ix2520 : xnor2 port map ( Y=>nx2519, A0=>nx1140, A1=>nx1238);
   ix1141 : oai32 port map ( Y=>nx1140, A0=>nx1567, A1=>nx1589, A2=>nx2349, 
      B0=>nx2523, B1=>nx2345);
   ix2524 : inv01 port map ( Y=>nx2523, A=>nx984);
   ix1239 : xnor2 port map ( Y=>nx1238, A0=>nx2527, A1=>nx1236);
   ix2528 : nand02 port map ( Y=>nx2527, A0=>nx3749, A1=>nx3705);
   ix1237 : xnor2 port map ( Y=>nx1236, A0=>nx1148, A1=>nx2533);
   ix1149 : oai32 port map ( Y=>nx1148, A0=>nx1855, A1=>nx1629, A2=>nx2357, 
      B0=>nx2351, B1=>nx2353);
   ix2534 : xnor2 port map ( Y=>nx2533, A0=>nx2535, A1=>nx2537);
   ix2536 : nand02 port map ( Y=>nx2535, A0=>nx3753, A1=>nx3701);
   ix2538 : xnor2 port map ( Y=>nx2537, A0=>nx2539, A1=>nx2541);
   ix2540 : aoi32 port map ( Y=>nx2539, A0=>nx3763, A1=>nx3697, A2=>nx1060, 
      B0=>nx1000, B1=>nx1062);
   ix2542 : xnor2 port map ( Y=>nx2541, A0=>nx2543, A1=>nx2545);
   ix2544 : nand02 port map ( Y=>nx2543, A0=>nx3757, A1=>nx3697);
   ix2546 : xnor2 port map ( Y=>nx2545, A0=>nx1164, A1=>nx1226);
   ix1165 : oai32 port map ( Y=>nx1164, A0=>nx1731, A1=>nx1703, A2=>nx2375, 
      B0=>nx2549, B1=>nx2371);
   ix2550 : inv01 port map ( Y=>nx2549, A=>nx1008);
   ix1227 : xnor2 port map ( Y=>nx1226, A0=>nx2553, A1=>nx1224);
   ix2554 : nand02 port map ( Y=>nx2553, A0=>nx3763, A1=>nx3693);
   ix1225 : xnor2 port map ( Y=>nx1224, A0=>nx1172, A1=>nx2559);
   ix1173 : oai32 port map ( Y=>nx1172, A0=>nx1579, A1=>nx1825, A2=>nx2383, 
      B0=>nx2377, B1=>nx2379);
   ix2560 : xnor2 port map ( Y=>nx2559, A0=>nx2561, A1=>nx2563);
   ix2562 : nand02 port map ( Y=>nx2561, A0=>nx3765, A1=>nx3689);
   ix2564 : xnor2 port map ( Y=>nx2563, A0=>nx2565, A1=>nx2567);
   ix2566 : aoi32 port map ( Y=>nx2565, A0=>nx3775, A1=>nx3685, A2=>nx1048, 
      B0=>nx1024, B1=>nx1050);
   ix2568 : xnor2 port map ( Y=>nx2567, A0=>nx2569, A1=>nx2571);
   ix2570 : nand02 port map ( Y=>nx2569, A0=>nx3769, A1=>nx3685);
   ix2572 : xnor2 port map ( Y=>nx2571, A0=>nx1188, A1=>nx1214);
   ix1189 : oai32 port map ( Y=>nx1188, A0=>nx1587, A1=>nx2165, A2=>nx2407, 
      B0=>nx2575, B1=>nx2403);
   ix2580 : inv01 port map ( Y=>nx2579, A=>A(13));
   ix1215 : xnor2 port map ( Y=>nx1214, A0=>nx2585, A1=>nx1212);
   ix2586 : nand02 port map ( Y=>nx2585, A0=>nx3775, A1=>nx3681);
   ix1213 : xnor2 port map ( Y=>nx1212, A0=>nx1196, A1=>nx2591);
   ix1197 : oai33 port map ( Y=>nx1196, A0=>nx1627, A1=>nx2391, A2=>nx2411, 
      B0=>nx1631, B1=>nx2579, B2=>nx2415);
   ix2592 : xnor2 port map ( Y=>nx2591, A0=>nx2593, A1=>nx2595);
   ix2594 : nand02 port map ( Y=>nx2593, A0=>nx3777, A1=>nx3677);
   ix2596 : xnor2 port map ( Y=>nx2595, A0=>nx2597, A1=>nx2599);
   ix2598 : nand02 port map ( Y=>nx2597, A0=>nx3781, A1=>nx3673);
   ix2600 : xnor2 port map ( Y=>nx2599, A0=>nx2601, A1=>nx2603);
   ix2602 : nand02 port map ( Y=>nx2601, A0=>nx3785, A1=>nx3669);
   ix2604 : nand02 port map ( Y=>nx2603, A0=>nx3665, A1=>nx3789);
   ix2879 : nor02ii port map ( Y=>Product(1), A0=>nx2607, A1=>nx2447);
   ix2608 : aoi22 port map ( Y=>nx2607, A0=>nx3723, A1=>nx3789, B0=>nx3787, 
      B1=>nx3727);
   ix2869 : xor2 port map ( Y=>Product(2), A0=>nx2447, A1=>nx2451);
   ix2863 : xor2 port map ( Y=>Product(3), A0=>nx14, A1=>nx36);
   ix2857 : xor2 port map ( Y=>Product(4), A0=>nx2443, A1=>nx2461);
   ix2851 : xnor2 port map ( Y=>Product(5), A0=>nx74, A1=>nx2439);
   ix2845 : xor2 port map ( Y=>Product(6), A0=>nx122, A1=>nx180);
   ix2839 : xor2 port map ( Y=>Product(7), A0=>nx2435, A1=>nx2465);
   ix2833 : xnor2 port map ( Y=>Product(8), A0=>nx254, A1=>nx2431);
   ix2827 : xor2 port map ( Y=>Product(9), A0=>nx338, A1=>nx432);
   ix2821 : xor2 port map ( Y=>Product(10), A0=>nx2427, A1=>nx2469);
   ix2815 : xnor2 port map ( Y=>Product(11), A0=>nx542, A1=>nx2423);
   ix2809 : xor2 port map ( Y=>Product(12), A0=>nx662, A1=>nx792);
   ix2803 : xor2 port map ( Y=>Product(13), A0=>nx2419, A1=>nx2473);
   ix2797 : xnor2 port map ( Y=>Product(14), A0=>nx938, A1=>nx1551);
   ix2785 : xor2 port map ( Y=>Product(16), A0=>nx2637, A1=>nx2639);
   ix2638 : nand02 port map ( Y=>nx2637, A0=>nx1094, A1=>nx1260);
   ix2640 : xnor2 port map ( Y=>nx2639, A0=>nx1268, A1=>nx1438);
   ix1269 : oai32 port map ( Y=>nx1268, A0=>nx2643, A1=>nx2195, A2=>nx2485, 
      B0=>nx2645, B1=>nx2481);
   ix2644 : inv01 port map ( Y=>nx2643, A=>B(15));
   ix2646 : inv01 port map ( Y=>nx2645, A=>nx1100);
   ix1439 : xnor2 port map ( Y=>nx1438, A0=>nx1274, A1=>nx2651);
   ix1275 : oai32 port map ( Y=>nx1274, A0=>nx2479, A1=>nx1561, A2=>nx2493, 
      B0=>nx2487, B1=>nx2489);
   ix2652 : xnor2 port map ( Y=>nx2651, A0=>nx2653, A1=>nx2655);
   ix2654 : nand02 port map ( Y=>nx2653, A0=>nx3729, A1=>nx3723);
   ix2656 : xnor2 port map ( Y=>nx2655, A0=>nx2657, A1=>nx2659);
   ix2658 : aoi32 port map ( Y=>nx2657, A0=>nx3737, A1=>nx3719, A2=>nx1248, 
      B0=>nx1116, B1=>nx1250);
   ix2660 : xnor2 port map ( Y=>nx2659, A0=>nx2661, A1=>nx2663);
   ix2662 : nand02 port map ( Y=>nx2661, A0=>nx3733, A1=>nx3719);
   ix2664 : xnor2 port map ( Y=>nx2663, A0=>nx1290, A1=>nx1428);
   ix1291 : oai32 port map ( Y=>nx1290, A0=>nx2193, A1=>nx1733, A2=>nx2511, 
      B0=>nx2667, B1=>nx2507);
   ix2668 : inv01 port map ( Y=>nx2667, A=>nx1124);
   ix1429 : xnor2 port map ( Y=>nx1428, A0=>nx2671, A1=>nx1426);
   ix2672 : nand02 port map ( Y=>nx2671, A0=>nx3737, A1=>nx3715);
   ix1427 : xnor2 port map ( Y=>nx1426, A0=>nx1298, A1=>nx2677);
   ix1299 : oai32 port map ( Y=>nx1298, A0=>nx1559, A1=>nx1581, A2=>nx2519, 
      B0=>nx2513, B1=>nx2515);
   ix2678 : xnor2 port map ( Y=>nx2677, A0=>nx2679, A1=>nx2681);
   ix2680 : nand02 port map ( Y=>nx2679, A0=>nx3741, A1=>nx3711);
   ix2682 : xnor2 port map ( Y=>nx2681, A0=>nx2683, A1=>nx2685);
   ix2684 : aoi32 port map ( Y=>nx2683, A0=>nx3749, A1=>nx3705, A2=>nx1236, 
      B0=>nx1140, B1=>nx1238);
   ix2686 : xnor2 port map ( Y=>nx2685, A0=>nx2687, A1=>nx2689);
   ix2688 : nand02 port map ( Y=>nx2687, A0=>nx3745, A1=>nx3705);
   ix2690 : xnor2 port map ( Y=>nx2689, A0=>nx1314, A1=>nx1416);
   ix1315 : oai32 port map ( Y=>nx1314, A0=>nx1567, A1=>nx1629, A2=>nx2537, 
      B0=>nx2693, B1=>nx2533);
   ix2694 : inv01 port map ( Y=>nx2693, A=>nx1148);
   ix1417 : xnor2 port map ( Y=>nx1416, A0=>nx2697, A1=>nx1414);
   ix2698 : nand02 port map ( Y=>nx2697, A0=>nx3749, A1=>nx3701);
   ix1415 : xnor2 port map ( Y=>nx1414, A0=>nx1322, A1=>nx2703);
   ix1323 : oai32 port map ( Y=>nx1322, A0=>nx1855, A1=>nx1605, A2=>nx2545, 
      B0=>nx2539, B1=>nx2541);
   ix2704 : xnor2 port map ( Y=>nx2703, A0=>nx2705, A1=>nx2707);
   ix2706 : nand02 port map ( Y=>nx2705, A0=>nx3753, A1=>nx3697);
   ix2708 : xnor2 port map ( Y=>nx2707, A0=>nx2709, A1=>nx2711);
   ix2710 : aoi32 port map ( Y=>nx2709, A0=>nx3763, A1=>nx3693, A2=>nx1224, 
      B0=>nx1164, B1=>nx1226);
   ix2712 : xnor2 port map ( Y=>nx2711, A0=>nx2713, A1=>nx2715);
   ix2714 : nand02 port map ( Y=>nx2713, A0=>nx3757, A1=>nx3693);
   ix2716 : xnor2 port map ( Y=>nx2715, A0=>nx1338, A1=>nx1404);
   ix1339 : oai32 port map ( Y=>nx1338, A0=>nx1731, A1=>nx1825, A2=>nx2563, 
      B0=>nx2719, B1=>nx2559);
   ix2720 : inv01 port map ( Y=>nx2719, A=>nx1172);
   ix1405 : xnor2 port map ( Y=>nx1404, A0=>nx2723, A1=>nx1402);
   ix2724 : nand02 port map ( Y=>nx2723, A0=>nx3763, A1=>nx3689);
   ix1403 : xnor2 port map ( Y=>nx1402, A0=>nx1346, A1=>nx2729);
   ix1347 : oai32 port map ( Y=>nx1346, A0=>nx1579, A1=>nx1979, A2=>nx2571, 
      B0=>nx2565, B1=>nx2567);
   ix2730 : xnor2 port map ( Y=>nx2729, A0=>nx2731, A1=>nx2733);
   ix2732 : nand02 port map ( Y=>nx2731, A0=>nx3765, A1=>nx3685);
   ix2734 : xnor2 port map ( Y=>nx2733, A0=>nx2735, A1=>nx2737);
   ix2736 : aoi32 port map ( Y=>nx2735, A0=>nx3775, A1=>nx3681, A2=>nx1212, 
      B0=>nx1188, B1=>nx1214);
   ix2738 : xnor2 port map ( Y=>nx2737, A0=>nx2739, A1=>nx2741);
   ix2740 : nand02 port map ( Y=>nx2739, A0=>nx3769, A1=>nx3681);
   ix2742 : xnor2 port map ( Y=>nx2741, A0=>nx1362, A1=>nx1392);
   ix1363 : oai32 port map ( Y=>nx1362, A0=>nx1587, A1=>nx2391, A2=>nx2595, 
      B0=>nx2745, B1=>nx2591);
   ix2750 : inv01 port map ( Y=>nx2749, A=>A(14));
   ix1393 : xnor2 port map ( Y=>nx1392, A0=>nx2755, A1=>nx1390);
   ix2756 : nand02 port map ( Y=>nx2755, A0=>nx3775, A1=>nx3677);
   ix1391 : xnor2 port map ( Y=>nx1390, A0=>nx1370, A1=>nx2763);
   ix1371 : oai33 port map ( Y=>nx1370, A0=>nx1627, A1=>nx2579, A2=>nx2599, 
      B0=>nx2601, B1=>nx2761, B2=>nx1607);
   ix2762 : inv01 port map ( Y=>nx2761, A=>A(15));
   ix2764 : xnor2 port map ( Y=>nx2763, A0=>nx2765, A1=>nx2767);
   ix2766 : nand02 port map ( Y=>nx2765, A0=>nx3777, A1=>nx3673);
   ix2768 : nand02 port map ( Y=>nx2767, A0=>nx2769, A1=>nx1382);
   ix2770 : nand04 port map ( Y=>nx2769, A0=>nx3781, A1=>nx3665, A2=>nx3787, 
      A3=>nx3669);
   ix2783 : xnor2 port map ( Y=>Product(17), A0=>nx2775, A1=>nx1604);
   ix2776 : aoi22 port map ( Y=>nx2775, A0=>nx1268, A1=>nx1438, B0=>nx1262, 
      B1=>nx1440);
   ix1605 : xnor2 port map ( Y=>nx1604, A0=>nx1452, A1=>nx2787);
   ix1453 : oai32 port map ( Y=>nx1452, A0=>nx2643, A1=>nx1561, A2=>nx2655, 
      B0=>nx2785, B1=>nx2651);
   ix2786 : inv01 port map ( Y=>nx2785, A=>nx1274);
   ix2788 : xnor2 port map ( Y=>nx2787, A0=>nx1458, A1=>nx1600);
   ix1459 : oai32 port map ( Y=>nx1458, A0=>nx2479, A1=>nx1569, A2=>nx2663, 
      B0=>nx2657, B1=>nx2659);
   ix1601 : xnor2 port map ( Y=>nx1600, A0=>nx2793, A1=>nx1598);
   ix2794 : nand02 port map ( Y=>nx2793, A0=>nx3729, A1=>nx3719);
   ix1599 : xnor2 port map ( Y=>nx1598, A0=>nx2797, A1=>nx1596);
   ix2798 : aoi32 port map ( Y=>nx2797, A0=>nx3737, A1=>nx3715, A2=>nx1426, 
      B0=>nx1290, B1=>nx1428);
   ix1597 : xnor2 port map ( Y=>nx1596, A0=>nx2801, A1=>nx1594);
   ix2802 : nand02 port map ( Y=>nx2801, A0=>nx3733, A1=>nx3715);
   ix1595 : xnor2 port map ( Y=>nx1594, A0=>nx1474, A1=>nx2809);
   ix1475 : oai32 port map ( Y=>nx1474, A0=>nx2193, A1=>nx1581, A2=>nx2681, 
      B0=>nx2807, B1=>nx2677);
   ix2808 : inv01 port map ( Y=>nx2807, A=>nx1298);
   ix2810 : xnor2 port map ( Y=>nx2809, A0=>nx2811, A1=>nx2813);
   ix2812 : nand02 port map ( Y=>nx2811, A0=>nx3737, A1=>nx3711);
   ix2814 : xnor2 port map ( Y=>nx2813, A0=>nx1482, A1=>nx1588);
   ix1483 : oai32 port map ( Y=>nx1482, A0=>nx1559, A1=>nx1589, A2=>nx2689, 
      B0=>nx2683, B1=>nx2685);
   ix1589 : xnor2 port map ( Y=>nx1588, A0=>nx2819, A1=>nx1586);
   ix2820 : nand02 port map ( Y=>nx2819, A0=>nx3741, A1=>nx3707);
   ix1587 : xnor2 port map ( Y=>nx1586, A0=>nx2823, A1=>nx1584);
   ix2824 : aoi32 port map ( Y=>nx2823, A0=>nx3749, A1=>nx3701, A2=>nx1414, 
      B0=>nx1314, B1=>nx1416);
   ix1585 : xnor2 port map ( Y=>nx1584, A0=>nx2827, A1=>nx1582);
   ix2828 : nand02 port map ( Y=>nx2827, A0=>nx3745, A1=>nx3701);
   ix1583 : xnor2 port map ( Y=>nx1582, A0=>nx1498, A1=>nx2835);
   ix1499 : oai32 port map ( Y=>nx1498, A0=>nx1567, A1=>nx1605, A2=>nx2707, 
      B0=>nx2833, B1=>nx2703);
   ix2834 : inv01 port map ( Y=>nx2833, A=>nx1322);
   ix2836 : xnor2 port map ( Y=>nx2835, A0=>nx2837, A1=>nx2839);
   ix2838 : nand02 port map ( Y=>nx2837, A0=>nx3749, A1=>nx3697);
   ix2840 : xnor2 port map ( Y=>nx2839, A0=>nx1506, A1=>nx1576);
   ix1507 : oai32 port map ( Y=>nx1506, A0=>nx1855, A1=>nx1703, A2=>nx2715, 
      B0=>nx2709, B1=>nx2711);
   ix1577 : xnor2 port map ( Y=>nx1576, A0=>nx2845, A1=>nx1574);
   ix2846 : nand02 port map ( Y=>nx2845, A0=>nx3753, A1=>nx3693);
   ix1575 : xnor2 port map ( Y=>nx1574, A0=>nx2849, A1=>nx1572);
   ix2850 : aoi32 port map ( Y=>nx2849, A0=>nx3763, A1=>nx3689, A2=>nx1402, 
      B0=>nx1338, B1=>nx1404);
   ix1573 : xnor2 port map ( Y=>nx1572, A0=>nx2853, A1=>nx1570);
   ix2854 : nand02 port map ( Y=>nx2853, A0=>nx3757, A1=>nx3689);
   ix1571 : xnor2 port map ( Y=>nx1570, A0=>nx1522, A1=>nx2861);
   ix1523 : oai32 port map ( Y=>nx1522, A0=>nx1731, A1=>nx1979, A2=>nx2733, 
      B0=>nx2859, B1=>nx2729);
   ix2860 : inv01 port map ( Y=>nx2859, A=>nx1346);
   ix2862 : xnor2 port map ( Y=>nx2861, A0=>nx2863, A1=>nx2865);
   ix2864 : nand02 port map ( Y=>nx2863, A0=>nx3763, A1=>nx3685);
   ix2866 : xnor2 port map ( Y=>nx2865, A0=>nx1530, A1=>nx1564);
   ix1531 : oai32 port map ( Y=>nx1530, A0=>nx1579, A1=>nx2165, A2=>nx2741, 
      B0=>nx2735, B1=>nx2737);
   ix1565 : xnor2 port map ( Y=>nx1564, A0=>nx2871, A1=>nx1562);
   ix2872 : nand02 port map ( Y=>nx2871, A0=>nx3765, A1=>nx3681);
   ix1563 : xnor2 port map ( Y=>nx1562, A0=>nx2875, A1=>nx1560);
   ix2876 : aoi32 port map ( Y=>nx2875, A0=>nx3775, A1=>nx3677, A2=>nx1390, 
      B0=>nx1362, B1=>nx1392);
   ix1561 : xnor2 port map ( Y=>nx1560, A0=>nx2879, A1=>nx1558);
   ix2880 : nand02 port map ( Y=>nx2879, A0=>nx3769, A1=>nx3677);
   ix1559 : xnor2 port map ( Y=>nx1558, A0=>nx1546, A1=>nx2887);
   ix1547 : oai32 port map ( Y=>nx1546, A0=>nx1587, A1=>nx2579, A2=>nx2767, 
      B0=>nx2883, B1=>nx2763);
   ix2888 : xnor2 port map ( Y=>nx2887, A0=>nx2889, A1=>nx2891);
   ix2890 : nand02 port map ( Y=>nx2889, A0=>nx3775, A1=>nx3673);
   ix2892 : xnor2 port map ( Y=>nx2891, A0=>nx2769, A1=>nx2893);
   ix2894 : xnor2 port map ( Y=>nx2893, A0=>nx2895, A1=>nx2897);
   ix2896 : nand02 port map ( Y=>nx2895, A0=>nx3777, A1=>nx3669);
   ix2898 : nand02 port map ( Y=>nx2897, A0=>nx3783, A1=>nx3665);
   ix2781 : xnor2 port map ( Y=>Product(18), A0=>nx2900, A1=>nx1764);
   ix2901 : aoi22 port map ( Y=>nx2900, A0=>nx1452, A1=>nx1602, B0=>nx1446, 
      B1=>nx1604);
   ix1765 : xnor2 port map ( Y=>nx1764, A0=>nx2907, A1=>nx1762);
   ix2908 : aoi32 port map ( Y=>nx2907, A0=>nx3729, A1=>nx3719, A2=>nx1598, 
      B0=>nx1458, B1=>nx1600);
   ix1763 : xnor2 port map ( Y=>nx1762, A0=>nx2910, A1=>nx1760);
   ix2911 : aoi32 port map ( Y=>nx2910, A0=>nx3733, A1=>nx3715, A2=>nx1594, 
      B0=>nx1466, B1=>nx1596);
   ix1761 : xnor2 port map ( Y=>nx1760, A0=>nx2914, A1=>nx1758);
   ix2915 : nand02 port map ( Y=>nx2914, A0=>nx3729, A1=>nx3715);
   ix1759 : xnor2 port map ( Y=>nx1758, A0=>nx1630, A1=>nx2924);
   ix1631 : oai32 port map ( Y=>nx1630, A0=>nx2918, A1=>nx1581, A2=>nx2813, 
      B0=>nx2920, B1=>nx2809);
   ix2919 : inv01 port map ( Y=>nx2918, A=>B(13));
   ix2925 : xnor2 port map ( Y=>nx2924, A0=>nx2926, A1=>nx2928);
   ix2927 : nand02 port map ( Y=>nx2926, A0=>nx3733, A1=>nx3711);
   ix2929 : xnor2 port map ( Y=>nx2928, A0=>nx2930, A1=>nx2932);
   ix2931 : aoi32 port map ( Y=>nx2930, A0=>nx3741, A1=>nx3707, A2=>nx1586, 
      B0=>nx1482, B1=>nx1588);
   ix2933 : xnor2 port map ( Y=>nx2932, A0=>nx2934, A1=>nx2936);
   ix2935 : nand02 port map ( Y=>nx2934, A0=>nx3737, A1=>nx3707);
   ix2937 : xnor2 port map ( Y=>nx2936, A0=>nx2938, A1=>nx2941);
   ix2939 : aoi32 port map ( Y=>nx2938, A0=>nx3745, A1=>nx3703, A2=>nx1582, 
      B0=>nx1490, B1=>nx1584);
   ix2942 : xnor2 port map ( Y=>nx2941, A0=>nx2943, A1=>nx2945);
   ix2944 : nand02 port map ( Y=>nx2943, A0=>nx3741, A1=>nx3703);
   ix2946 : xnor2 port map ( Y=>nx2945, A0=>nx1654, A1=>nx1744);
   ix1655 : oai32 port map ( Y=>nx1654, A0=>nx2948, A1=>nx1605, A2=>nx2839, 
      B0=>nx2950, B1=>nx2835);
   ix2949 : inv01 port map ( Y=>nx2948, A=>B(10));
   ix1745 : xnor2 port map ( Y=>nx1744, A0=>nx2955, A1=>nx1742);
   ix2956 : nand02 port map ( Y=>nx2955, A0=>nx3745, A1=>nx3697);
   ix1743 : xnor2 port map ( Y=>nx1742, A0=>nx2958, A1=>nx1740);
   ix2959 : aoi32 port map ( Y=>nx2958, A0=>nx3753, A1=>nx3693, A2=>nx1574, 
      B0=>nx1506, B1=>nx1576);
   ix1741 : xnor2 port map ( Y=>nx1740, A0=>nx2961, A1=>nx1738);
   ix2962 : nand02 port map ( Y=>nx2961, A0=>nx3751, A1=>nx3693);
   ix1739 : xnor2 port map ( Y=>nx1738, A0=>nx2964, A1=>nx1736);
   ix2965 : aoi32 port map ( Y=>nx2964, A0=>nx3757, A1=>nx3689, A2=>nx1570, 
      B0=>nx1514, B1=>nx1572);
   ix1737 : xnor2 port map ( Y=>nx1736, A0=>nx2968, A1=>nx1734);
   ix2969 : nand02 port map ( Y=>nx2968, A0=>nx3753, A1=>nx3689);
   ix1735 : xnor2 port map ( Y=>nx1734, A0=>nx1678, A1=>nx2978);
   ix1679 : oai32 port map ( Y=>nx1678, A0=>nx2972, A1=>nx1979, A2=>nx2865, 
      B0=>nx2974, B1=>nx2861);
   ix2973 : inv01 port map ( Y=>nx2972, A=>B(7));
   ix2979 : xnor2 port map ( Y=>nx2978, A0=>nx2980, A1=>nx2982);
   ix2981 : nand02 port map ( Y=>nx2980, A0=>nx3757, A1=>nx3685);
   ix2983 : xnor2 port map ( Y=>nx2982, A0=>nx2984, A1=>nx2986);
   ix2985 : aoi32 port map ( Y=>nx2984, A0=>nx3765, A1=>nx3681, A2=>nx1562, 
      B0=>nx1530, B1=>nx1564);
   ix2987 : xnor2 port map ( Y=>nx2986, A0=>nx2988, A1=>nx2990);
   ix2989 : nand02 port map ( Y=>nx2988, A0=>nx3763, A1=>nx3681);
   ix2991 : xnor2 port map ( Y=>nx2990, A0=>nx2992, A1=>nx2995);
   ix2993 : aoi32 port map ( Y=>nx2992, A0=>nx3769, A1=>nx3677, A2=>nx1558, 
      B0=>nx1538, B1=>nx1560);
   ix2996 : xnor2 port map ( Y=>nx2995, A0=>nx2997, A1=>nx2999);
   ix2998 : nand02 port map ( Y=>nx2997, A0=>nx3765, A1=>nx3677);
   ix3000 : xnor2 port map ( Y=>nx2999, A0=>nx1702, A1=>nx1720);
   ix1703 : oai32 port map ( Y=>nx1702, A0=>nx3002, A1=>nx2579, A2=>nx2891, 
      B0=>nx3004, B1=>nx2887);
   ix3003 : inv01 port map ( Y=>nx3002, A=>B(4));
   ix3008 : aoi22 port map ( Y=>nx3007, A0=>nx3787, A1=>nx3665, B0=>nx3783, 
      B1=>nx3669);
   ix1721 : xnor2 port map ( Y=>nx1720, A0=>nx3011, A1=>nx1718);
   ix3012 : nand02 port map ( Y=>nx3011, A0=>nx3769, A1=>nx3673);
   ix1719 : xnor2 port map ( Y=>nx1718, A0=>nx1710, A1=>nx3015);
   ix1711 : aoi21 port map ( Y=>nx1710, A0=>nx2895, A1=>nx2601, B0=>nx2897);
   ix3016 : xnor2 port map ( Y=>nx3015, A0=>nx3017, A1=>nx3019);
   ix3018 : nand02 port map ( Y=>nx3017, A0=>nx3775, A1=>nx3669);
   ix3020 : nand02 port map ( Y=>nx3019, A0=>nx3779, A1=>nx3665);
   ix2779 : xor2 port map ( Y=>Product(19), A0=>nx1770, A1=>nx1912);
   ix1771 : oai22 port map ( Y=>nx1770, A0=>nx2900, A1=>nx3023, B0=>nx2907, 
      B1=>nx3025);
   ix1913 : xnor2 port map ( Y=>nx1912, A0=>nx3028, A1=>nx1910);
   ix3029 : aoi32 port map ( Y=>nx3028, A0=>nx3729, A1=>nx3715, A2=>nx1758, 
      B0=>nx1622, B1=>nx1760);
   ix1911 : xnor2 port map ( Y=>nx1910, A0=>nx1782, A1=>nx3037);
   ix1783 : oai32 port map ( Y=>nx1782, A0=>nx2479, A1=>nx1581, A2=>nx2928, 
      B0=>nx3033, B1=>nx2924);
   ix3038 : xnor2 port map ( Y=>nx3037, A0=>nx3039, A1=>nx3041);
   ix3040 : nand02 port map ( Y=>nx3039, A0=>nx3729, A1=>nx3711);
   ix3042 : xnor2 port map ( Y=>nx3041, A0=>nx1790, A1=>nx1904);
   ix1791 : oai32 port map ( Y=>nx1790, A0=>nx2918, A1=>nx1589, A2=>nx2936, 
      B0=>nx2930, B1=>nx2932);
   ix1905 : xnor2 port map ( Y=>nx1904, A0=>nx3045, A1=>nx1902);
   ix3046 : nand02 port map ( Y=>nx3045, A0=>nx3733, A1=>nx3707);
   ix1903 : xnor2 port map ( Y=>nx1902, A0=>nx1798, A1=>nx3049);
   ix1799 : oai32 port map ( Y=>nx1798, A0=>nx2193, A1=>nx1629, A2=>nx2945, 
      B0=>nx2938, B1=>nx2941);
   ix3050 : xnor2 port map ( Y=>nx3049, A0=>nx3051, A1=>nx3053);
   ix3052 : nand02 port map ( Y=>nx3051, A0=>nx3737, A1=>nx3703);
   ix3054 : xnor2 port map ( Y=>nx3053, A0=>nx3055, A1=>nx3057);
   ix3056 : aoi32 port map ( Y=>nx3055, A0=>nx3745, A1=>nx3697, A2=>nx1742, 
      B0=>nx1654, B1=>nx1744);
   ix3058 : xnor2 port map ( Y=>nx3057, A0=>nx3059, A1=>nx3061);
   ix3060 : nand02 port map ( Y=>nx3059, A0=>nx3741, A1=>nx3699);
   ix3062 : xnor2 port map ( Y=>nx3061, A0=>nx3063, A1=>nx3066);
   ix3064 : aoi32 port map ( Y=>nx3063, A0=>nx3751, A1=>nx3693, A2=>nx1738, 
      B0=>nx1662, B1=>nx1740);
   ix3067 : xnor2 port map ( Y=>nx3066, A0=>nx3068, A1=>nx3070);
   ix3069 : nand02 port map ( Y=>nx3068, A0=>nx3745, A1=>nx3695);
   ix3071 : xnor2 port map ( Y=>nx3070, A0=>nx3072, A1=>nx3075);
   ix3073 : aoi32 port map ( Y=>nx3072, A0=>nx3753, A1=>nx3689, A2=>nx1734, 
      B0=>nx1670, B1=>nx1736);
   ix3076 : xnor2 port map ( Y=>nx3075, A0=>nx3077, A1=>nx3079);
   ix3078 : nand02 port map ( Y=>nx3077, A0=>nx3751, A1=>nx3689);
   ix3080 : xnor2 port map ( Y=>nx3079, A0=>nx1830, A1=>nx1884);
   ix1831 : oai32 port map ( Y=>nx1830, A0=>nx1855, A1=>nx1979, A2=>nx2982, 
      B0=>nx3082, B1=>nx2978);
   ix1885 : xnor2 port map ( Y=>nx1884, A0=>nx3087, A1=>nx1882);
   ix3088 : nand02 port map ( Y=>nx3087, A0=>nx3753, A1=>nx3685);
   ix1883 : xnor2 port map ( Y=>nx1882, A0=>nx1838, A1=>nx3091);
   ix1839 : oai32 port map ( Y=>nx1838, A0=>nx2972, A1=>nx2165, A2=>nx2990, 
      B0=>nx2984, B1=>nx2986);
   ix3092 : xnor2 port map ( Y=>nx3091, A0=>nx3093, A1=>nx3095);
   ix3094 : nand02 port map ( Y=>nx3093, A0=>nx3757, A1=>nx3681);
   ix3096 : xnor2 port map ( Y=>nx3095, A0=>nx1846, A1=>nx1876);
   ix1847 : oai32 port map ( Y=>nx1846, A0=>nx1731, A1=>nx2391, A2=>nx2999, 
      B0=>nx2992, B1=>nx2995);
   ix1877 : xnor2 port map ( Y=>nx1876, A0=>nx3099, A1=>nx1874);
   ix3100 : nand02 port map ( Y=>nx3099, A0=>nx3763, A1=>nx3677);
   ix1875 : xnor2 port map ( Y=>nx1874, A0=>nx3102, A1=>nx1872);
   ix3103 : aoi32 port map ( Y=>nx3102, A0=>nx3771, A1=>nx3673, A2=>nx1718, 
      B0=>nx1702, B1=>nx1720);
   ix1873 : xnor2 port map ( Y=>nx1872, A0=>nx3105, A1=>nx1870);
   ix3106 : nand02 port map ( Y=>nx3105, A0=>nx3765, A1=>nx3673);
   ix1871 : xnor2 port map ( Y=>nx1870, A0=>nx1862, A1=>nx3111);
   ix1863 : oai32 port map ( Y=>nx1862, A0=>nx3002, A1=>nx2749, A2=>nx3019, 
      B0=>nx3109, B1=>nx3015);
   ix3112 : xnor2 port map ( Y=>nx3111, A0=>nx3113, A1=>nx3115);
   ix3114 : nand02 port map ( Y=>nx3113, A0=>nx3771, A1=>nx3669);
   ix3116 : nand02 port map ( Y=>nx3115, A0=>nx3775, A1=>nx3665);
   ix2777 : xnor2 port map ( Y=>Product(20), A0=>nx3118, A1=>nx2048);
   ix3119 : aoi22 port map ( Y=>nx3118, A0=>nx1776, A1=>nx1910, B0=>nx1770, 
      B1=>nx1912);
   ix2049 : xnor2 port map ( Y=>nx2048, A0=>nx1924, A1=>nx3127);
   ix1925 : oai32 port map ( Y=>nx1924, A0=>nx2643, A1=>nx1581, A2=>nx3041, 
      B0=>nx3123, B1=>nx3037);
   ix3128 : xnor2 port map ( Y=>nx3127, A0=>nx3129, A1=>nx3131);
   ix3130 : aoi32 port map ( Y=>nx3129, A0=>nx3733, A1=>nx3707, A2=>nx1902, 
      B0=>nx1790, B1=>nx1904);
   ix3132 : xnor2 port map ( Y=>nx3131, A0=>nx3133, A1=>nx3135);
   ix3134 : nand02 port map ( Y=>nx3133, A0=>nx3729, A1=>nx3707);
   ix3136 : xnor2 port map ( Y=>nx3135, A0=>nx1938, A1=>nx2040);
   ix1939 : oai32 port map ( Y=>nx1938, A0=>nx2918, A1=>nx1629, A2=>nx3053, 
      B0=>nx3138, B1=>nx3049);
   ix3139 : inv01 port map ( Y=>nx3138, A=>nx1798);
   ix2041 : xnor2 port map ( Y=>nx2040, A0=>nx3141, A1=>nx2038);
   ix3142 : nand02 port map ( Y=>nx3141, A0=>nx3733, A1=>nx3703);
   ix2039 : xnor2 port map ( Y=>nx2038, A0=>nx1946, A1=>nx3145);
   ix1947 : oai32 port map ( Y=>nx1946, A0=>nx2193, A1=>nx1605, A2=>nx3061, 
      B0=>nx3055, B1=>nx3057);
   ix3146 : xnor2 port map ( Y=>nx3145, A0=>nx3147, A1=>nx3149);
   ix3148 : nand02 port map ( Y=>nx3147, A0=>nx3737, A1=>nx3699);
   ix3150 : xnor2 port map ( Y=>nx3149, A0=>nx1954, A1=>nx2032);
   ix1955 : oai32 port map ( Y=>nx1954, A0=>nx1559, A1=>nx1703, A2=>nx3070, 
      B0=>nx3063, B1=>nx3066);
   ix2033 : xnor2 port map ( Y=>nx2032, A0=>nx3153, A1=>nx2030);
   ix3154 : nand02 port map ( Y=>nx3153, A0=>nx3741, A1=>nx3695);
   ix2031 : xnor2 port map ( Y=>nx2030, A0=>nx1962, A1=>nx3157);
   ix1963 : oai32 port map ( Y=>nx1962, A0=>nx2948, A1=>nx1825, A2=>nx3079, 
      B0=>nx3072, B1=>nx3075);
   ix3158 : xnor2 port map ( Y=>nx3157, A0=>nx3159, A1=>nx3161);
   ix3160 : nand02 port map ( Y=>nx3159, A0=>nx3745, A1=>nx3691);
   ix3162 : xnor2 port map ( Y=>nx3161, A0=>nx3163, A1=>nx3165);
   ix3164 : aoi32 port map ( Y=>nx3163, A0=>nx3753, A1=>nx3685, A2=>nx1882, 
      B0=>nx1830, B1=>nx1884);
   ix3166 : xnor2 port map ( Y=>nx3165, A0=>nx3167, A1=>nx3169);
   ix3168 : nand02 port map ( Y=>nx3167, A0=>nx3751, A1=>nx3685);
   ix3170 : xnor2 port map ( Y=>nx3169, A0=>nx1978, A1=>nx2020);
   ix1979 : oai32 port map ( Y=>nx1978, A0=>nx1855, A1=>nx2165, A2=>nx3095, 
      B0=>nx3172, B1=>nx3091);
   ix3173 : inv01 port map ( Y=>nx3172, A=>nx1838);
   ix2021 : xnor2 port map ( Y=>nx2020, A0=>nx3175, A1=>nx2018);
   ix3176 : nand02 port map ( Y=>nx3175, A0=>nx3753, A1=>nx3681);
   ix2019 : xnor2 port map ( Y=>nx2018, A0=>nx3178, A1=>nx2016);
   ix3179 : aoi32 port map ( Y=>nx3178, A0=>nx3763, A1=>nx3677, A2=>nx1874, 
      B0=>nx1846, B1=>nx1876);
   ix2017 : xnor2 port map ( Y=>nx2016, A0=>nx3181, A1=>nx2014);
   ix3182 : nand02 port map ( Y=>nx3181, A0=>nx3757, A1=>nx3677);
   ix2015 : xnor2 port map ( Y=>nx2014, A0=>nx3184, A1=>nx2012);
   ix3185 : aoi32 port map ( Y=>nx3184, A0=>nx3767, A1=>nx3673, A2=>nx1870, 
      B0=>nx1854, B1=>nx1872);
   ix2013 : xnor2 port map ( Y=>nx2012, A0=>nx3188, A1=>nx2010);
   ix3189 : nand02 port map ( Y=>nx3188, A0=>nx3763, A1=>nx3673);
   ix2011 : xnor2 port map ( Y=>nx2010, A0=>nx2002, A1=>nx3196);
   ix2003 : oai32 port map ( Y=>nx2002, A0=>nx1579, A1=>nx2749, A2=>nx3115, 
      B0=>nx3192, B1=>nx3111);
   ix3197 : xnor2 port map ( Y=>nx3196, A0=>nx3198, A1=>nx3200);
   ix3199 : nand02 port map ( Y=>nx3198, A0=>nx3767, A1=>nx3669);
   ix3201 : nand02 port map ( Y=>nx3200, A0=>nx3771, A1=>nx3665);
   ix2775 : xor2 port map ( Y=>Product(21), A0=>nx2054, A1=>nx2172);
   ix2055 : oai22 port map ( Y=>nx2054, A0=>nx3118, A1=>nx3204, B0=>nx3206, 
      B1=>nx3127);
   ix2173 : xnor2 port map ( Y=>nx2172, A0=>nx2060, A1=>nx3212);
   ix2061 : oai32 port map ( Y=>nx2060, A0=>nx2643, A1=>nx1589, A2=>nx3135, 
      B0=>nx3129, B1=>nx3131);
   ix3213 : xnor2 port map ( Y=>nx3212, A0=>nx3214, A1=>nx3216);
   ix3215 : aoi32 port map ( Y=>nx3214, A0=>nx3733, A1=>nx3703, A2=>nx2038, 
      B0=>nx1938, B1=>nx2040);
   ix3217 : xnor2 port map ( Y=>nx3216, A0=>nx3218, A1=>nx3220);
   ix3219 : nand02 port map ( Y=>nx3218, A0=>nx3729, A1=>nx3703);
   ix3221 : xnor2 port map ( Y=>nx3220, A0=>nx2074, A1=>nx2164);
   ix2075 : oai32 port map ( Y=>nx2074, A0=>nx2918, A1=>nx1605, A2=>nx3149, 
      B0=>nx3223, B1=>nx3145);
   ix3224 : inv01 port map ( Y=>nx3223, A=>nx1946);
   ix2165 : xnor2 port map ( Y=>nx2164, A0=>nx3226, A1=>nx2162);
   ix3227 : nand02 port map ( Y=>nx3226, A0=>nx3733, A1=>nx3699);
   ix2163 : xnor2 port map ( Y=>nx2162, A0=>nx3229, A1=>nx2160);
   ix3230 : aoi32 port map ( Y=>nx3229, A0=>nx3741, A1=>nx3695, A2=>nx2030, 
      B0=>nx1954, B1=>nx2032);
   ix2161 : xnor2 port map ( Y=>nx2160, A0=>nx3232, A1=>nx2158);
   ix3233 : nand02 port map ( Y=>nx3232, A0=>nx3737, A1=>nx3695);
   ix2159 : xnor2 port map ( Y=>nx2158, A0=>nx2090, A1=>nx3238);
   ix2091 : oai32 port map ( Y=>nx2090, A0=>nx1559, A1=>nx1825, A2=>nx3161, 
      B0=>nx3236, B1=>nx3157);
   ix3237 : inv01 port map ( Y=>nx3236, A=>nx1962);
   ix3239 : xnor2 port map ( Y=>nx3238, A0=>nx3240, A1=>nx3242);
   ix3241 : nand02 port map ( Y=>nx3240, A0=>nx3741, A1=>nx3691);
   ix3243 : xnor2 port map ( Y=>nx3242, A0=>nx2098, A1=>nx2152);
   ix2099 : oai32 port map ( Y=>nx2098, A0=>nx2948, A1=>nx1979, A2=>nx3169, 
      B0=>nx3163, B1=>nx3165);
   ix2153 : xnor2 port map ( Y=>nx2152, A0=>nx3246, A1=>nx2150);
   ix3247 : nand02 port map ( Y=>nx3246, A0=>nx3745, A1=>nx3685);
   ix2151 : xnor2 port map ( Y=>nx2150, A0=>nx3249, A1=>nx2148);
   ix3250 : aoi32 port map ( Y=>nx3249, A0=>nx3755, A1=>nx3681, A2=>nx2018, 
      B0=>nx1978, B1=>nx2020);
   ix2149 : xnor2 port map ( Y=>nx2148, A0=>nx3252, A1=>nx2146);
   ix3253 : nand02 port map ( Y=>nx3252, A0=>nx3751, A1=>nx3681);
   ix2147 : xnor2 port map ( Y=>nx2146, A0=>nx3255, A1=>nx2144);
   ix3256 : aoi32 port map ( Y=>nx3255, A0=>nx3757, A1=>nx3677, A2=>nx2014, 
      B0=>nx1986, B1=>nx2016);
   ix2145 : xnor2 port map ( Y=>nx2144, A0=>nx3259, A1=>nx2142);
   ix3260 : nand02 port map ( Y=>nx3259, A0=>nx3755, A1=>nx3677);
   ix2143 : xnor2 port map ( Y=>nx2142, A0=>nx3262, A1=>nx2140);
   ix3263 : aoi32 port map ( Y=>nx3262, A0=>nx3763, A1=>nx3673, A2=>nx2010, 
      B0=>nx1994, B1=>nx2012);
   ix2141 : xnor2 port map ( Y=>nx2140, A0=>nx3266, A1=>nx2138);
   ix3267 : nand02 port map ( Y=>nx3266, A0=>nx3759, A1=>nx3673);
   ix2139 : xnor2 port map ( Y=>nx2138, A0=>nx2130, A1=>nx3274);
   ix2131 : oai32 port map ( Y=>nx2130, A0=>nx1731, A1=>nx2749, A2=>nx3200, 
      B0=>nx3270, B1=>nx3196);
   ix3275 : xnor2 port map ( Y=>nx3274, A0=>nx3276, A1=>nx3278);
   ix3277 : nand02 port map ( Y=>nx3276, A0=>nx3763, A1=>nx3669);
   ix3279 : nand02 port map ( Y=>nx3278, A0=>nx3767, A1=>nx3665);
   ix2773 : xnor2 port map ( Y=>Product(22), A0=>nx3281, A1=>nx2284);
   ix3282 : aoi22 port map ( Y=>nx3281, A0=>nx2060, A1=>nx2170, B0=>nx2054, 
      B1=>nx2172);
   ix2285 : xnor2 port map ( Y=>nx2284, A0=>nx2184, A1=>nx3286);
   ix2185 : oai32 port map ( Y=>nx2184, A0=>nx2643, A1=>nx1629, A2=>nx3220, 
      B0=>nx3214, B1=>nx3216);
   ix3287 : xnor2 port map ( Y=>nx3286, A0=>nx3288, A1=>nx3290);
   ix3289 : aoi32 port map ( Y=>nx3288, A0=>nx3733, A1=>nx3699, A2=>nx2162, 
      B0=>nx2074, B1=>nx2164);
   ix3291 : xnor2 port map ( Y=>nx3290, A0=>nx3292, A1=>nx3294);
   ix3293 : nand02 port map ( Y=>nx3292, A0=>nx3729, A1=>nx3699);
   ix3295 : xnor2 port map ( Y=>nx3294, A0=>nx3296, A1=>nx3299);
   ix3297 : aoi32 port map ( Y=>nx3296, A0=>nx3737, A1=>nx3695, A2=>nx2158, 
      B0=>nx2082, B1=>nx2160);
   ix3300 : xnor2 port map ( Y=>nx3299, A0=>nx3301, A1=>nx3303);
   ix3302 : nand02 port map ( Y=>nx3301, A0=>nx3733, A1=>nx3695);
   ix3304 : xnor2 port map ( Y=>nx3303, A0=>nx2206, A1=>nx2272);
   ix2207 : oai32 port map ( Y=>nx2206, A0=>nx2193, A1=>nx1825, A2=>nx3242, 
      B0=>nx3306, B1=>nx3238);
   ix2273 : xnor2 port map ( Y=>nx2272, A0=>nx3311, A1=>nx2270);
   ix3312 : nand02 port map ( Y=>nx3311, A0=>nx3737, A1=>nx3691);
   ix2271 : xnor2 port map ( Y=>nx2270, A0=>nx3314, A1=>nx2268);
   ix3315 : aoi32 port map ( Y=>nx3314, A0=>nx3745, A1=>nx3685, A2=>nx2150, 
      B0=>nx2098, B1=>nx2152);
   ix2269 : xnor2 port map ( Y=>nx2268, A0=>nx3317, A1=>nx2266);
   ix3318 : nand02 port map ( Y=>nx3317, A0=>nx3741, A1=>nx3687);
   ix2267 : xnor2 port map ( Y=>nx2266, A0=>nx3320, A1=>nx2264);
   ix3321 : aoi32 port map ( Y=>nx3320, A0=>nx3751, A1=>nx3681, A2=>nx2146, 
      B0=>nx2106, B1=>nx2148);
   ix2265 : xnor2 port map ( Y=>nx2264, A0=>nx3324, A1=>nx2262);
   ix3325 : nand02 port map ( Y=>nx3324, A0=>nx3745, A1=>nx3683);
   ix2263 : xnor2 port map ( Y=>nx2262, A0=>nx3327, A1=>nx2260);
   ix3328 : aoi32 port map ( Y=>nx3327, A0=>nx3755, A1=>nx3677, A2=>nx2142, 
      B0=>nx2114, B1=>nx2144);
   ix2261 : xnor2 port map ( Y=>nx2260, A0=>nx3331, A1=>nx2258);
   ix3332 : nand02 port map ( Y=>nx3331, A0=>nx3751, A1=>nx3679);
   ix2259 : xnor2 port map ( Y=>nx2258, A0=>nx3334, A1=>nx2256);
   ix3335 : aoi32 port map ( Y=>nx3334, A0=>nx3759, A1=>nx3673, A2=>nx2138, 
      B0=>nx2122, B1=>nx2140);
   ix2257 : xnor2 port map ( Y=>nx2256, A0=>nx3338, A1=>nx2254);
   ix3339 : nand02 port map ( Y=>nx3338, A0=>nx3755, A1=>nx3673);
   ix2255 : xnor2 port map ( Y=>nx2254, A0=>nx2246, A1=>nx3346);
   ix2247 : oai32 port map ( Y=>nx2246, A0=>nx2972, A1=>nx2749, A2=>nx3278, 
      B0=>nx3342, B1=>nx3274);
   ix3347 : xnor2 port map ( Y=>nx3346, A0=>nx3348, A1=>nx3350);
   ix3349 : nand02 port map ( Y=>nx3348, A0=>nx3759, A1=>nx3669);
   ix3351 : nand02 port map ( Y=>nx3350, A0=>nx3763, A1=>nx3665);
   ix2771 : xor2 port map ( Y=>Product(23), A0=>nx2290, A1=>nx2384);
   ix2291 : oai22 port map ( Y=>nx2290, A0=>nx3281, A1=>nx3354, B0=>nx3356, 
      B1=>nx3286);
   ix3357 : inv01 port map ( Y=>nx3356, A=>nx2184);
   ix2385 : xnor2 port map ( Y=>nx2384, A0=>nx2296, A1=>nx3360);
   ix2297 : oai32 port map ( Y=>nx2296, A0=>nx2643, A1=>nx1605, A2=>nx3294, 
      B0=>nx3288, B1=>nx3290);
   ix3361 : xnor2 port map ( Y=>nx3360, A0=>nx2302, A1=>nx2380);
   ix2303 : oai32 port map ( Y=>nx2302, A0=>nx2479, A1=>nx1703, A2=>nx3303, 
      B0=>nx3296, B1=>nx3299);
   ix2381 : xnor2 port map ( Y=>nx2380, A0=>nx3364, A1=>nx2378);
   ix3365 : nand02 port map ( Y=>nx3364, A0=>nx3729, A1=>nx3695);
   ix2379 : xnor2 port map ( Y=>nx2378, A0=>nx3367, A1=>nx2376);
   ix3368 : aoi32 port map ( Y=>nx3367, A0=>nx3739, A1=>nx3691, A2=>nx2270, 
      B0=>nx2206, B1=>nx2272);
   ix2377 : xnor2 port map ( Y=>nx2376, A0=>nx3370, A1=>nx2374);
   ix3371 : nand02 port map ( Y=>nx3370, A0=>nx3733, A1=>nx3691);
   ix2375 : xnor2 port map ( Y=>nx2374, A0=>nx3373, A1=>nx2372);
   ix3374 : aoi32 port map ( Y=>nx3373, A0=>nx3741, A1=>nx3687, A2=>nx2266, 
      B0=>nx2214, B1=>nx2268);
   ix2373 : xnor2 port map ( Y=>nx2372, A0=>nx3377, A1=>nx2370);
   ix3378 : nand02 port map ( Y=>nx3377, A0=>nx3739, A1=>nx3687);
   ix2371 : xnor2 port map ( Y=>nx2370, A0=>nx3380, A1=>nx2368);
   ix3381 : aoi32 port map ( Y=>nx3380, A0=>nx3747, A1=>nx3683, A2=>nx2262, 
      B0=>nx2222, B1=>nx2264);
   ix2369 : xnor2 port map ( Y=>nx2368, A0=>nx3384, A1=>nx2366);
   ix3385 : nand02 port map ( Y=>nx3384, A0=>nx3741, A1=>nx3683);
   ix2367 : xnor2 port map ( Y=>nx2366, A0=>nx3387, A1=>nx2364);
   ix3388 : aoi32 port map ( Y=>nx3387, A0=>nx3751, A1=>nx3679, A2=>nx2258, 
      B0=>nx2230, B1=>nx2260);
   ix2365 : xnor2 port map ( Y=>nx2364, A0=>nx3391, A1=>nx2362);
   ix3392 : nand02 port map ( Y=>nx3391, A0=>nx3747, A1=>nx3679);
   ix2363 : xnor2 port map ( Y=>nx2362, A0=>nx3394, A1=>nx2360);
   ix3395 : aoi32 port map ( Y=>nx3394, A0=>nx3755, A1=>nx3673, A2=>nx2254, 
      B0=>nx2238, B1=>nx2256);
   ix2361 : xnor2 port map ( Y=>nx2360, A0=>nx3398, A1=>nx2358);
   ix3399 : nand02 port map ( Y=>nx3398, A0=>nx3751, A1=>nx3675);
   ix2359 : xnor2 port map ( Y=>nx2358, A0=>nx2350, A1=>nx3406);
   ix2351 : oai32 port map ( Y=>nx2350, A0=>nx1855, A1=>nx2749, A2=>nx3350, 
      B0=>nx3402, B1=>nx3346);
   ix3407 : xnor2 port map ( Y=>nx3406, A0=>nx3408, A1=>nx3410);
   ix3409 : nand02 port map ( Y=>nx3408, A0=>nx3755, A1=>nx3669);
   ix3411 : nand02 port map ( Y=>nx3410, A0=>nx3759, A1=>nx3665);
   ix2769 : xnor2 port map ( Y=>Product(24), A0=>nx3413, A1=>nx2472);
   ix3414 : aoi22 port map ( Y=>nx3413, A0=>nx2296, A1=>nx2382, B0=>nx2290, 
      B1=>nx2384);
   ix2473 : xnor2 port map ( Y=>nx2472, A0=>nx3417, A1=>nx2470);
   ix3418 : aoi32 port map ( Y=>nx3417, A0=>nx3729, A1=>nx3695, A2=>nx2378, 
      B0=>nx2302, B1=>nx2380);
   ix2471 : xnor2 port map ( Y=>nx2470, A0=>nx3420, A1=>nx2468);
   ix3421 : aoi32 port map ( Y=>nx3420, A0=>nx3733, A1=>nx3691, A2=>nx2374, 
      B0=>nx2310, B1=>nx2376);
   ix2469 : xnor2 port map ( Y=>nx2468, A0=>nx3424, A1=>nx2466);
   ix3425 : nand02 port map ( Y=>nx3424, A0=>nx3729, A1=>nx3691);
   ix2467 : xnor2 port map ( Y=>nx2466, A0=>nx3427, A1=>nx2464);
   ix3428 : aoi32 port map ( Y=>nx3427, A0=>nx3739, A1=>nx3687, A2=>nx2370, 
      B0=>nx2318, B1=>nx2372);
   ix2465 : xnor2 port map ( Y=>nx2464, A0=>nx3431, A1=>nx2462);
   ix3432 : nand02 port map ( Y=>nx3431, A0=>nx3735, A1=>nx3687);
   ix2463 : xnor2 port map ( Y=>nx2462, A0=>nx3434, A1=>nx2460);
   ix3435 : aoi32 port map ( Y=>nx3434, A0=>nx3743, A1=>nx3683, A2=>nx2366, 
      B0=>nx2326, B1=>nx2368);
   ix2461 : xnor2 port map ( Y=>nx2460, A0=>nx3438, A1=>nx2458);
   ix3439 : nand02 port map ( Y=>nx3438, A0=>nx3739, A1=>nx3683);
   ix2459 : xnor2 port map ( Y=>nx2458, A0=>nx3441, A1=>nx2456);
   ix3442 : aoi32 port map ( Y=>nx3441, A0=>nx3747, A1=>nx3679, A2=>nx2362, 
      B0=>nx2334, B1=>nx2364);
   ix2457 : xnor2 port map ( Y=>nx2456, A0=>nx3445, A1=>nx2454);
   ix3446 : nand02 port map ( Y=>nx3445, A0=>nx3743, A1=>nx3679);
   ix2455 : xnor2 port map ( Y=>nx2454, A0=>nx3448, A1=>nx2452);
   ix3449 : aoi32 port map ( Y=>nx3448, A0=>nx3751, A1=>nx3675, A2=>nx2358, 
      B0=>nx2342, B1=>nx2360);
   ix2453 : xnor2 port map ( Y=>nx2452, A0=>nx3452, A1=>nx2450);
   ix3453 : nand02 port map ( Y=>nx3452, A0=>nx3747, A1=>nx3675);
   ix2451 : xnor2 port map ( Y=>nx2450, A0=>nx2442, A1=>nx3460);
   ix2443 : oai32 port map ( Y=>nx2442, A0=>nx1567, A1=>nx2749, A2=>nx3410, 
      B0=>nx3456, B1=>nx3406);
   ix3461 : xnor2 port map ( Y=>nx3460, A0=>nx3462, A1=>nx3464);
   ix3463 : nand02 port map ( Y=>nx3462, A0=>nx3751, A1=>nx3669);
   ix3465 : nand02 port map ( Y=>nx3464, A0=>nx3755, A1=>nx3665);
   ix2767 : xor2 port map ( Y=>Product(25), A0=>nx2478, A1=>nx2548);
   ix2479 : oai22 port map ( Y=>nx2478, A0=>nx3413, A1=>nx3468, B0=>nx3417, 
      B1=>nx3470);
   ix2549 : xnor2 port map ( Y=>nx2548, A0=>nx3473, A1=>nx2546);
   ix3474 : aoi32 port map ( Y=>nx3473, A0=>nx3729, A1=>nx3691, A2=>nx2466, 
      B0=>nx2402, B1=>nx2468);
   ix2547 : xnor2 port map ( Y=>nx2546, A0=>nx3477, A1=>nx2544);
   ix3478 : aoi32 port map ( Y=>nx3477, A0=>nx3735, A1=>nx3687, A2=>nx2462, 
      B0=>nx2410, B1=>nx2464);
   ix2545 : xnor2 port map ( Y=>nx2544, A0=>nx3481, A1=>nx2542);
   ix3482 : nand02 port map ( Y=>nx3481, A0=>nx3729, A1=>nx3687);
   ix2543 : xnor2 port map ( Y=>nx2542, A0=>nx3484, A1=>nx2540);
   ix3485 : aoi32 port map ( Y=>nx3484, A0=>nx3739, A1=>nx3683, A2=>nx2458, 
      B0=>nx2418, B1=>nx2460);
   ix2541 : xnor2 port map ( Y=>nx2540, A0=>nx3488, A1=>nx2538);
   ix3489 : nand02 port map ( Y=>nx3488, A0=>nx3735, A1=>nx3683);
   ix2539 : xnor2 port map ( Y=>nx2538, A0=>nx3491, A1=>nx2536);
   ix3492 : aoi32 port map ( Y=>nx3491, A0=>nx3743, A1=>nx3679, A2=>nx2454, 
      B0=>nx2426, B1=>nx2456);
   ix2537 : xnor2 port map ( Y=>nx2536, A0=>nx3495, A1=>nx2534);
   ix3496 : nand02 port map ( Y=>nx3495, A0=>nx3739, A1=>nx3679);
   ix2535 : xnor2 port map ( Y=>nx2534, A0=>nx3498, A1=>nx2532);
   ix3499 : aoi32 port map ( Y=>nx3498, A0=>nx3747, A1=>nx3675, A2=>nx2450, 
      B0=>nx2434, B1=>nx2452);
   ix2533 : xnor2 port map ( Y=>nx2532, A0=>nx3502, A1=>nx2530);
   ix3503 : nand02 port map ( Y=>nx3502, A0=>nx3743, A1=>nx3675);
   ix2531 : xnor2 port map ( Y=>nx2530, A0=>nx2522, A1=>nx3510);
   ix2523 : oai32 port map ( Y=>nx2522, A0=>nx2948, A1=>nx2749, A2=>nx3464, 
      B0=>nx3506, B1=>nx3460);
   ix3511 : xnor2 port map ( Y=>nx3510, A0=>nx3512, A1=>nx3514);
   ix3513 : nand02 port map ( Y=>nx3512, A0=>nx3747, A1=>nx3669);
   ix3515 : nand02 port map ( Y=>nx3514, A0=>nx3751, A1=>nx3665);
   ix2765 : xnor2 port map ( Y=>Product(26), A0=>nx3517, A1=>nx2612);
   ix3518 : aoi22 port map ( Y=>nx3517, A0=>nx2484, A1=>nx2546, B0=>nx2478, 
      B1=>nx2548);
   ix2613 : xnor2 port map ( Y=>nx2612, A0=>nx3521, A1=>nx2610);
   ix3522 : aoi32 port map ( Y=>nx3521, A0=>nx3731, A1=>nx3687, A2=>nx2542, 
      B0=>nx2490, B1=>nx2544);
   ix2611 : xnor2 port map ( Y=>nx2610, A0=>nx3525, A1=>nx2608);
   ix3526 : aoi32 port map ( Y=>nx3525, A0=>nx3735, A1=>nx3683, A2=>nx2538, 
      B0=>nx2498, B1=>nx2540);
   ix2609 : xnor2 port map ( Y=>nx2608, A0=>nx3529, A1=>nx2606);
   ix3530 : nand02 port map ( Y=>nx3529, A0=>nx3731, A1=>nx3683);
   ix2607 : xnor2 port map ( Y=>nx2606, A0=>nx3532, A1=>nx2604);
   ix3533 : aoi32 port map ( Y=>nx3532, A0=>nx3739, A1=>nx3679, A2=>nx2534, 
      B0=>nx2506, B1=>nx2536);
   ix2605 : xnor2 port map ( Y=>nx2604, A0=>nx3536, A1=>nx2602);
   ix3537 : nand02 port map ( Y=>nx3536, A0=>nx3735, A1=>nx3679);
   ix2603 : xnor2 port map ( Y=>nx2602, A0=>nx3539, A1=>nx2600);
   ix3540 : aoi32 port map ( Y=>nx3539, A0=>nx3743, A1=>nx3675, A2=>nx2530, 
      B0=>nx2514, B1=>nx2532);
   ix2601 : xnor2 port map ( Y=>nx2600, A0=>nx3543, A1=>nx2598);
   ix3544 : nand02 port map ( Y=>nx3543, A0=>nx3739, A1=>nx3675);
   ix2599 : xnor2 port map ( Y=>nx2598, A0=>nx2590, A1=>nx3551);
   ix2591 : oai32 port map ( Y=>nx2590, A0=>nx1559, A1=>nx2749, A2=>nx3514, 
      B0=>nx3547, B1=>nx3510);
   ix3552 : xnor2 port map ( Y=>nx3551, A0=>nx3553, A1=>nx3555);
   ix3554 : nand02 port map ( Y=>nx3553, A0=>nx3743, A1=>nx3669);
   ix3556 : nand02 port map ( Y=>nx3555, A0=>nx3747, A1=>nx3665);
   ix2763 : xor2 port map ( Y=>Product(27), A0=>nx2618, A1=>nx2664);
   ix2619 : oai22 port map ( Y=>nx2618, A0=>nx3517, A1=>nx3559, B0=>nx3521, 
      B1=>nx3561);
   ix2665 : xnor2 port map ( Y=>nx2664, A0=>nx3564, A1=>nx2662);
   ix3565 : aoi32 port map ( Y=>nx3564, A0=>nx3731, A1=>nx3683, A2=>nx2606, 
      B0=>nx2566, B1=>nx2608);
   ix2663 : xnor2 port map ( Y=>nx2662, A0=>nx3568, A1=>nx2660);
   ix3569 : aoi32 port map ( Y=>nx3568, A0=>nx3735, A1=>nx3679, A2=>nx2602, 
      B0=>nx2574, B1=>nx2604);
   ix2661 : xnor2 port map ( Y=>nx2660, A0=>nx3572, A1=>nx2658);
   ix3573 : nand02 port map ( Y=>nx3572, A0=>nx3731, A1=>nx3679);
   ix2659 : xnor2 port map ( Y=>nx2658, A0=>nx3575, A1=>nx2656);
   ix3576 : aoi32 port map ( Y=>nx3575, A0=>nx3739, A1=>nx3675, A2=>nx2598, 
      B0=>nx2582, B1=>nx2600);
   ix2657 : xnor2 port map ( Y=>nx2656, A0=>nx3579, A1=>nx2654);
   ix3580 : nand02 port map ( Y=>nx3579, A0=>nx3735, A1=>nx3675);
   ix2655 : xnor2 port map ( Y=>nx2654, A0=>nx2646, A1=>nx3587);
   ix2647 : oai32 port map ( Y=>nx2646, A0=>nx2193, A1=>nx2749, A2=>nx3555, 
      B0=>nx3583, B1=>nx3551);
   ix3588 : xnor2 port map ( Y=>nx3587, A0=>nx3589, A1=>nx3591);
   ix3590 : nand02 port map ( Y=>nx3589, A0=>nx3739, A1=>nx3669);
   ix3592 : nand02 port map ( Y=>nx3591, A0=>nx3743, A1=>nx3665);
   ix2761 : xnor2 port map ( Y=>Product(28), A0=>nx3594, A1=>nx2704);
   ix3595 : aoi22 port map ( Y=>nx3594, A0=>nx2624, A1=>nx2662, B0=>nx2618, 
      B1=>nx2664);
   ix2705 : xnor2 port map ( Y=>nx2704, A0=>nx3598, A1=>nx2702);
   ix3599 : aoi32 port map ( Y=>nx3598, A0=>nx3731, A1=>nx3679, A2=>nx2658, 
      B0=>nx2630, B1=>nx2660);
   ix2703 : xnor2 port map ( Y=>nx2702, A0=>nx3602, A1=>nx2700);
   ix3603 : aoi32 port map ( Y=>nx3602, A0=>nx3735, A1=>nx3675, A2=>nx2654, 
      B0=>nx2638, B1=>nx2656);
   ix2701 : xnor2 port map ( Y=>nx2700, A0=>nx3606, A1=>nx2698);
   ix3607 : nand02 port map ( Y=>nx3606, A0=>nx3731, A1=>nx3675);
   ix2699 : xnor2 port map ( Y=>nx2698, A0=>nx2690, A1=>nx3614);
   ix2691 : oai32 port map ( Y=>nx2690, A0=>nx2918, A1=>nx2749, A2=>nx3591, 
      B0=>nx3610, B1=>nx3587);
   ix3615 : xnor2 port map ( Y=>nx3614, A0=>nx3616, A1=>nx3618);
   ix3617 : nand02 port map ( Y=>nx3616, A0=>nx3735, A1=>nx3671);
   ix3619 : nand02 port map ( Y=>nx3618, A0=>nx3739, A1=>nx3665);
   ix2759 : xor2 port map ( Y=>Product(29), A0=>nx2710, A1=>nx2732);
   ix2711 : oai22 port map ( Y=>nx2710, A0=>nx3594, A1=>nx3622, B0=>nx3598, 
      B1=>nx3624);
   ix2733 : xnor2 port map ( Y=>nx2732, A0=>nx3627, A1=>nx2730);
   ix3628 : aoi32 port map ( Y=>nx3627, A0=>nx3731, A1=>nx3675, A2=>nx2698, 
      B0=>nx2682, B1=>nx2700);
   ix2731 : xnor2 port map ( Y=>nx2730, A0=>nx2722, A1=>nx3636);
   ix2723 : oai32 port map ( Y=>nx2722, A0=>nx2479, A1=>nx2749, A2=>nx3618, 
      B0=>nx3632, B1=>nx3614);
   ix3637 : xnor2 port map ( Y=>nx3636, A0=>nx3638, A1=>nx3640);
   ix3639 : nand02 port map ( Y=>nx3638, A0=>nx3731, A1=>nx3671);
   ix3641 : nand02 port map ( Y=>nx3640, A0=>nx3735, A1=>nx3667);
   ix2751 : xnor2 port map ( Y=>Product(30), A0=>nx3643, A1=>nx2748);
   ix3644 : aoi22 port map ( Y=>nx3643, A0=>nx2716, A1=>nx2730, B0=>nx2710, 
      B1=>nx2732);
   ix2749 : xnor2 port map ( Y=>nx2748, A0=>nx2744, A1=>nx3652);
   ix2745 : oai32 port map ( Y=>nx2744, A0=>nx2643, A1=>nx2749, A2=>nx3640, 
      B0=>nx3648, B1=>nx3636);
   ix3653 : nand02 port map ( Y=>nx3652, A0=>nx3731, A1=>nx3667);
   ix2757 : ao32 port map ( Y=>Product(31), A0=>nx2744, A1=>nx3731, A2=>
      nx3667, B0=>nx2738, B1=>nx2748);
   ix2739 : inv01 port map ( Y=>nx2738, A=>nx3643);
   ix3649 : inv01 port map ( Y=>nx3648, A=>nx2722);
   ix2717 : inv01 port map ( Y=>nx2716, A=>nx3627);
   ix3623 : inv01 port map ( Y=>nx3622, A=>nx2704);
   ix3625 : inv01 port map ( Y=>nx3624, A=>nx2702);
   ix3633 : inv01 port map ( Y=>nx3632, A=>nx2690);
   ix2683 : inv01 port map ( Y=>nx2682, A=>nx3602);
   ix3611 : inv01 port map ( Y=>nx3610, A=>nx2646);
   ix2639 : inv01 port map ( Y=>nx2638, A=>nx3575);
   ix2631 : inv01 port map ( Y=>nx2630, A=>nx3568);
   ix2625 : inv01 port map ( Y=>nx2624, A=>nx3564);
   ix3560 : inv01 port map ( Y=>nx3559, A=>nx2612);
   ix3562 : inv01 port map ( Y=>nx3561, A=>nx2610);
   ix3584 : inv01 port map ( Y=>nx3583, A=>nx2590);
   ix2583 : inv01 port map ( Y=>nx2582, A=>nx3539);
   ix2575 : inv01 port map ( Y=>nx2574, A=>nx3532);
   ix2567 : inv01 port map ( Y=>nx2566, A=>nx3525);
   ix3548 : inv01 port map ( Y=>nx3547, A=>nx2522);
   ix2515 : inv01 port map ( Y=>nx2514, A=>nx3498);
   ix2507 : inv01 port map ( Y=>nx2506, A=>nx3491);
   ix2499 : inv01 port map ( Y=>nx2498, A=>nx3484);
   ix2491 : inv01 port map ( Y=>nx2490, A=>nx3477);
   ix2485 : inv01 port map ( Y=>nx2484, A=>nx3473);
   ix3469 : inv01 port map ( Y=>nx3468, A=>nx2472);
   ix3471 : inv01 port map ( Y=>nx3470, A=>nx2470);
   ix3507 : inv01 port map ( Y=>nx3506, A=>nx2442);
   ix2435 : inv01 port map ( Y=>nx2434, A=>nx3448);
   ix2427 : inv01 port map ( Y=>nx2426, A=>nx3441);
   ix2419 : inv01 port map ( Y=>nx2418, A=>nx3434);
   ix2411 : inv01 port map ( Y=>nx2410, A=>nx3427);
   ix2403 : inv01 port map ( Y=>nx2402, A=>nx3420);
   ix2383 : inv01 port map ( Y=>nx2382, A=>nx3360);
   ix3457 : inv01 port map ( Y=>nx3456, A=>nx2350);
   ix2343 : inv01 port map ( Y=>nx2342, A=>nx3394);
   ix2335 : inv01 port map ( Y=>nx2334, A=>nx3387);
   ix2327 : inv01 port map ( Y=>nx2326, A=>nx3380);
   ix2319 : inv01 port map ( Y=>nx2318, A=>nx3373);
   ix2311 : inv01 port map ( Y=>nx2310, A=>nx3367);
   ix3355 : inv01 port map ( Y=>nx3354, A=>nx2284);
   ix3403 : inv01 port map ( Y=>nx3402, A=>nx2246);
   ix2239 : inv01 port map ( Y=>nx2238, A=>nx3334);
   ix2231 : inv01 port map ( Y=>nx2230, A=>nx3327);
   ix2223 : inv01 port map ( Y=>nx2222, A=>nx3320);
   ix2215 : inv01 port map ( Y=>nx2214, A=>nx3314);
   ix2171 : inv01 port map ( Y=>nx2170, A=>nx3212);
   ix3343 : inv01 port map ( Y=>nx3342, A=>nx2130);
   ix2123 : inv01 port map ( Y=>nx2122, A=>nx3262);
   ix2115 : inv01 port map ( Y=>nx2114, A=>nx3255);
   ix2107 : inv01 port map ( Y=>nx2106, A=>nx3249);
   ix3307 : inv01 port map ( Y=>nx3306, A=>nx2090);
   ix2083 : inv01 port map ( Y=>nx2082, A=>nx3229);
   ix3205 : inv01 port map ( Y=>nx3204, A=>nx2048);
   ix3271 : inv01 port map ( Y=>nx3270, A=>nx2002);
   ix1995 : inv01 port map ( Y=>nx1994, A=>nx3184);
   ix1987 : inv01 port map ( Y=>nx1986, A=>nx3178);
   ix3207 : inv01 port map ( Y=>nx3206, A=>nx1924);
   ix3193 : inv01 port map ( Y=>nx3192, A=>nx1862);
   ix1855 : inv01 port map ( Y=>nx1854, A=>nx3102);
   ix3124 : inv01 port map ( Y=>nx3123, A=>nx1782);
   ix1777 : inv01 port map ( Y=>nx1776, A=>nx3028);
   ix3024 : inv01 port map ( Y=>nx3023, A=>nx1764);
   ix3026 : inv01 port map ( Y=>nx3025, A=>nx1762);
   ix3110 : inv01 port map ( Y=>nx3109, A=>nx1710);
   ix3083 : inv01 port map ( Y=>nx3082, A=>nx1678);
   ix1671 : inv01 port map ( Y=>nx1670, A=>nx2964);
   ix1663 : inv01 port map ( Y=>nx1662, A=>nx2958);
   ix3034 : inv01 port map ( Y=>nx3033, A=>nx1630);
   ix1623 : inv01 port map ( Y=>nx1622, A=>nx2910);
   ix1603 : inv01 port map ( Y=>nx1602, A=>nx2787);
   ix3005 : inv01 port map ( Y=>nx3004, A=>nx1546);
   ix1539 : inv01 port map ( Y=>nx1538, A=>nx2875);
   ix2975 : inv01 port map ( Y=>nx2974, A=>nx1522);
   ix1515 : inv01 port map ( Y=>nx1514, A=>nx2849);
   ix2951 : inv01 port map ( Y=>nx2950, A=>nx1498);
   ix1491 : inv01 port map ( Y=>nx1490, A=>nx2823);
   ix2921 : inv01 port map ( Y=>nx2920, A=>nx1474);
   ix1467 : inv01 port map ( Y=>nx1466, A=>nx2797);
   ix1447 : inv01 port map ( Y=>nx1446, A=>nx2775);
   ix1441 : inv01 port map ( Y=>nx1440, A=>nx2639);
   ix1383 : inv01 port map ( Y=>nx1382, A=>nx3007);
   ix2884 : inv01 port map ( Y=>nx2883, A=>nx1370);
   ix1263 : inv01 port map ( Y=>nx1262, A=>nx2637);
   ix2746 : inv01 port map ( Y=>nx2745, A=>nx1196);
   ix2576 : inv01 port map ( Y=>nx2575, A=>nx1032);
   ix2388 : inv01 port map ( Y=>nx2387, A=>nx880);
   ix2162 : inv01 port map ( Y=>nx2161, A=>nx740);
   ix1976 : inv01 port map ( Y=>nx1975, A=>nx612);
   ix1822 : inv01 port map ( Y=>nx1821, A=>nx496);
   ix1700 : inv01 port map ( Y=>nx1699, A=>nx392);
   ix1602 : inv01 port map ( Y=>nx1601, A=>nx300);
   ix1662 : inv01 port map ( Y=>nx1661, A=>nx220);
   ix1758 : inv01 port map ( Y=>nx1757, A=>nx152);
   ix1888 : inv01 port map ( Y=>nx1887, A=>nx96);
   ix2048 : inv01 port map ( Y=>nx2047, A=>nx52);
   ix2248 : inv01 port map ( Y=>nx2247, A=>nx20);
   ix3 : and02 port map ( Y=>Product_0_EXMPLR, A0=>nx3791, A1=>nx3727);
   ix3664 : inv01 port map ( Y=>nx3665, A=>nx2761);
   ix3666 : inv01 port map ( Y=>nx3667, A=>nx2761);
   ix3668 : inv01 port map ( Y=>nx3669, A=>nx2749);
   ix3670 : inv01 port map ( Y=>nx3671, A=>nx2749);
   ix3672 : inv01 port map ( Y=>nx3673, A=>nx2579);
   ix3674 : inv01 port map ( Y=>nx3675, A=>nx2579);
   ix3676 : inv01 port map ( Y=>nx3677, A=>nx2391);
   ix3678 : inv01 port map ( Y=>nx3679, A=>nx2391);
   ix3680 : inv01 port map ( Y=>nx3681, A=>nx2165);
   ix3682 : inv01 port map ( Y=>nx3683, A=>nx2165);
   ix3684 : inv01 port map ( Y=>nx3685, A=>nx1979);
   ix3686 : inv01 port map ( Y=>nx3687, A=>nx1979);
   ix3688 : inv01 port map ( Y=>nx3689, A=>nx1825);
   ix3690 : inv01 port map ( Y=>nx3691, A=>nx1825);
   ix3692 : inv01 port map ( Y=>nx3693, A=>nx1703);
   ix3694 : inv01 port map ( Y=>nx3695, A=>nx1703);
   ix3696 : inv01 port map ( Y=>nx3697, A=>nx1605);
   ix3698 : inv01 port map ( Y=>nx3699, A=>nx1605);
   ix3700 : inv01 port map ( Y=>nx3701, A=>nx1629);
   ix3702 : inv01 port map ( Y=>nx3703, A=>nx1629);
   ix3704 : inv01 port map ( Y=>nx3705, A=>nx1589);
   ix3706 : inv01 port map ( Y=>nx3707, A=>nx1589);
   ix3708 : inv01 port map ( Y=>nx3709, A=>nx1581);
   ix3710 : inv01 port map ( Y=>nx3711, A=>nx1581);
   ix3712 : inv01 port map ( Y=>nx3713, A=>nx1733);
   ix3714 : inv01 port map ( Y=>nx3715, A=>nx1733);
   ix3716 : inv01 port map ( Y=>nx3717, A=>nx1569);
   ix3718 : inv01 port map ( Y=>nx3719, A=>nx1569);
   ix3720 : inv01 port map ( Y=>nx3721, A=>nx1561);
   ix3722 : inv01 port map ( Y=>nx3723, A=>nx1561);
   ix3724 : inv01 port map ( Y=>nx3725, A=>nx2195);
   ix3726 : inv01 port map ( Y=>nx3727, A=>nx2195);
   ix3728 : inv01 port map ( Y=>nx3729, A=>nx2643);
   ix3730 : inv01 port map ( Y=>nx3731, A=>nx2643);
   ix3732 : inv01 port map ( Y=>nx3733, A=>nx2479);
   ix3734 : inv01 port map ( Y=>nx3735, A=>nx2479);
   ix3736 : inv01 port map ( Y=>nx3737, A=>nx2918);
   ix3738 : inv01 port map ( Y=>nx3739, A=>nx2918);
   ix3740 : inv01 port map ( Y=>nx3741, A=>nx2193);
   ix3742 : inv01 port map ( Y=>nx3743, A=>nx2193);
   ix3744 : inv01 port map ( Y=>nx3745, A=>nx1559);
   ix3746 : inv01 port map ( Y=>nx3747, A=>nx1559);
   ix3748 : inv01 port map ( Y=>nx3749, A=>nx2948);
   ix3750 : inv01 port map ( Y=>nx3751, A=>nx2948);
   ix3752 : inv01 port map ( Y=>nx3753, A=>nx1567);
   ix3754 : inv01 port map ( Y=>nx3755, A=>nx1567);
   ix3756 : inv01 port map ( Y=>nx3757, A=>nx1855);
   ix3758 : inv01 port map ( Y=>nx3759, A=>nx1855);
   ix3760 : inv01 port map ( Y=>nx3761, A=>nx2972);
   ix3762 : inv01 port map ( Y=>nx3763, A=>nx2972);
   ix3764 : inv01 port map ( Y=>nx3765, A=>nx1731);
   ix3766 : inv01 port map ( Y=>nx3767, A=>nx1731);
   ix3768 : inv01 port map ( Y=>nx3769, A=>nx1579);
   ix3770 : inv01 port map ( Y=>nx3771, A=>nx1579);
   ix3772 : inv01 port map ( Y=>nx3773, A=>nx3002);
   ix3774 : inv01 port map ( Y=>nx3775, A=>nx3002);
   ix3776 : inv01 port map ( Y=>nx3777, A=>nx1587);
   ix3778 : inv01 port map ( Y=>nx3779, A=>nx1587);
   ix3780 : inv01 port map ( Y=>nx3781, A=>nx1627);
   ix3782 : inv01 port map ( Y=>nx3783, A=>nx1627);
   ix3784 : inv01 port map ( Y=>nx3785, A=>nx1631);
   ix3786 : inv01 port map ( Y=>nx3787, A=>nx1631);
   ix3788 : inv01 port map ( Y=>nx3789, A=>nx1607);
   ix3790 : inv01 port map ( Y=>nx3791, A=>nx1607);
end structural ;

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity RCFA_32 is
   port (
      A : IN std_logic_vector (31 DOWNTO 0) ;
      B : IN std_logic_vector (31 DOWNTO 0) ;
      Cin : IN std_logic ;
      Sum : OUT std_logic_vector (31 DOWNTO 0) ;
      Cout : OUT std_logic) ;
end RCFA_32 ;

architecture structural of RCFA_32 is
   signal nx8, nx10, nx12, nx22, nx28, nx30, nx32, nx42, nx48, nx50, nx52, 
      nx62, nx68, nx70, nx72, nx82, nx88, nx90, nx92, nx102, nx108, nx110, 
      nx112, nx122, nx128, nx130, nx132, nx142, nx148, nx150, nx152, nx162, 
      nx168, nx170, nx172, nx182, nx188, nx190, nx192, nx202, nx208, nx210, 
      nx212, nx222, nx228, nx230, nx232, nx242, nx248, nx250, nx252, nx262, 
      nx268, nx270, nx272, nx282, nx288, nx290, nx292, nx302, nx308, nx310, 
      nx312, nx510, nx514, nx518, nx522, nx526, nx530, nx534, nx538, nx542, 
      nx546, nx550, nx554, nx558, nx562, nx566, nx571, nx573, nx575, nx577, 
      nx580, nx582, nx584, nx586, nx589, nx591, nx593, nx595, nx598, nx600, 
      nx602, nx604, nx607, nx609, nx611, nx613, nx616, nx618, nx620, nx622, 
      nx625, nx627, nx629, nx631, nx634, nx636, nx638, nx640, nx643, nx645, 
      nx647, nx649, nx652, nx654, nx656, nx658, nx661, nx663, nx665, nx667, 
      nx670, nx672, nx674, nx676, nx679, nx681, nx683, nx685, nx688, nx690, 
      nx692, nx694, nx697, nx699, nx701, nx703, nx706: std_logic ;

begin
   ix321 : ao22 port map ( Y=>Cout, A0=>A(31), A1=>nx310, B0=>nx308, B1=>
      nx312);
   ix309 : oai22 port map ( Y=>nx308, A0=>nx510, A1=>nx699, B0=>nx703, B1=>
      nx701);
   ix511 : aoi22 port map ( Y=>nx510, A0=>A(29), A1=>nx290, B0=>nx288, B1=>
      nx292);
   ix289 : oai22 port map ( Y=>nx288, A0=>nx514, A1=>nx690, B0=>nx694, B1=>
      nx692);
   ix515 : aoi22 port map ( Y=>nx514, A0=>A(27), A1=>nx270, B0=>nx268, B1=>
      nx272);
   ix269 : oai22 port map ( Y=>nx268, A0=>nx518, A1=>nx681, B0=>nx685, B1=>
      nx683);
   ix519 : aoi22 port map ( Y=>nx518, A0=>A(25), A1=>nx250, B0=>nx248, B1=>
      nx252);
   ix249 : oai22 port map ( Y=>nx248, A0=>nx522, A1=>nx672, B0=>nx676, B1=>
      nx674);
   ix523 : aoi22 port map ( Y=>nx522, A0=>A(23), A1=>nx230, B0=>nx228, B1=>
      nx232);
   ix229 : oai22 port map ( Y=>nx228, A0=>nx526, A1=>nx663, B0=>nx667, B1=>
      nx665);
   ix527 : aoi22 port map ( Y=>nx526, A0=>A(21), A1=>nx210, B0=>nx208, B1=>
      nx212);
   ix209 : oai22 port map ( Y=>nx208, A0=>nx530, A1=>nx654, B0=>nx658, B1=>
      nx656);
   ix531 : aoi22 port map ( Y=>nx530, A0=>A(19), A1=>nx190, B0=>nx188, B1=>
      nx192);
   ix189 : oai22 port map ( Y=>nx188, A0=>nx534, A1=>nx645, B0=>nx649, B1=>
      nx647);
   ix535 : aoi22 port map ( Y=>nx534, A0=>A(17), A1=>nx170, B0=>nx168, B1=>
      nx172);
   ix169 : oai22 port map ( Y=>nx168, A0=>nx538, A1=>nx636, B0=>nx640, B1=>
      nx638);
   ix539 : aoi22 port map ( Y=>nx538, A0=>A(15), A1=>nx150, B0=>nx148, B1=>
      nx152);
   ix149 : oai22 port map ( Y=>nx148, A0=>nx542, A1=>nx627, B0=>nx631, B1=>
      nx629);
   ix543 : aoi22 port map ( Y=>nx542, A0=>A(13), A1=>nx130, B0=>nx128, B1=>
      nx132);
   ix129 : oai22 port map ( Y=>nx128, A0=>nx546, A1=>nx618, B0=>nx622, B1=>
      nx620);
   ix547 : aoi22 port map ( Y=>nx546, A0=>A(11), A1=>nx110, B0=>nx108, B1=>
      nx112);
   ix109 : oai22 port map ( Y=>nx108, A0=>nx550, A1=>nx609, B0=>nx613, B1=>
      nx611);
   ix551 : aoi22 port map ( Y=>nx550, A0=>A(9), A1=>nx90, B0=>nx88, B1=>nx92
   );
   ix89 : oai22 port map ( Y=>nx88, A0=>nx554, A1=>nx600, B0=>nx604, B1=>
      nx602);
   ix555 : aoi22 port map ( Y=>nx554, A0=>A(7), A1=>nx70, B0=>nx68, B1=>nx72
   );
   ix69 : oai22 port map ( Y=>nx68, A0=>nx558, A1=>nx591, B0=>nx595, B1=>
      nx593);
   ix559 : aoi22 port map ( Y=>nx558, A0=>A(5), A1=>nx50, B0=>nx48, B1=>nx52
   );
   ix49 : oai22 port map ( Y=>nx48, A0=>nx562, A1=>nx582, B0=>nx586, B1=>
      nx584);
   ix563 : aoi22 port map ( Y=>nx562, A0=>A(3), A1=>nx30, B0=>nx28, B1=>nx32
   );
   ix29 : oai22 port map ( Y=>nx28, A0=>nx566, A1=>nx573, B0=>nx577, B1=>
      nx575);
   ix567 : aoi22 port map ( Y=>nx566, A0=>A(1), A1=>nx10, B0=>nx8, B1=>nx12
   );
   ix9 : mux21 port map ( Y=>nx8, A0=>Cin, A1=>A(0), S0=>B(0));
   ix13 : xnor2 port map ( Y=>nx12, A0=>A(1), A1=>nx571);
   ix572 : xnor2 port map ( Y=>nx571, A0=>B(1), A1=>Cin);
   ix576 : xnor2 port map ( Y=>nx575, A0=>B(2), A1=>Cin);
   ix578 : inv01 port map ( Y=>nx577, A=>A(2));
   ix33 : xnor2 port map ( Y=>nx32, A0=>A(3), A1=>nx580);
   ix581 : xnor2 port map ( Y=>nx580, A0=>B(3), A1=>Cin);
   ix585 : xnor2 port map ( Y=>nx584, A0=>B(4), A1=>Cin);
   ix587 : inv01 port map ( Y=>nx586, A=>A(4));
   ix53 : xnor2 port map ( Y=>nx52, A0=>A(5), A1=>nx589);
   ix590 : xnor2 port map ( Y=>nx589, A0=>B(5), A1=>Cin);
   ix594 : xnor2 port map ( Y=>nx593, A0=>B(6), A1=>Cin);
   ix596 : inv01 port map ( Y=>nx595, A=>A(6));
   ix73 : xnor2 port map ( Y=>nx72, A0=>A(7), A1=>nx598);
   ix599 : xnor2 port map ( Y=>nx598, A0=>B(7), A1=>Cin);
   ix603 : xnor2 port map ( Y=>nx602, A0=>B(8), A1=>Cin);
   ix605 : inv01 port map ( Y=>nx604, A=>A(8));
   ix93 : xnor2 port map ( Y=>nx92, A0=>A(9), A1=>nx607);
   ix608 : xnor2 port map ( Y=>nx607, A0=>B(9), A1=>Cin);
   ix612 : xnor2 port map ( Y=>nx611, A0=>B(10), A1=>Cin);
   ix614 : inv01 port map ( Y=>nx613, A=>A(10));
   ix113 : xnor2 port map ( Y=>nx112, A0=>A(11), A1=>nx616);
   ix617 : xnor2 port map ( Y=>nx616, A0=>B(11), A1=>Cin);
   ix621 : xnor2 port map ( Y=>nx620, A0=>B(12), A1=>Cin);
   ix623 : inv01 port map ( Y=>nx622, A=>A(12));
   ix133 : xnor2 port map ( Y=>nx132, A0=>A(13), A1=>nx625);
   ix626 : xnor2 port map ( Y=>nx625, A0=>B(13), A1=>Cin);
   ix630 : xnor2 port map ( Y=>nx629, A0=>B(14), A1=>Cin);
   ix632 : inv01 port map ( Y=>nx631, A=>A(14));
   ix153 : xnor2 port map ( Y=>nx152, A0=>A(15), A1=>nx634);
   ix635 : xnor2 port map ( Y=>nx634, A0=>B(15), A1=>Cin);
   ix639 : xnor2 port map ( Y=>nx638, A0=>B(16), A1=>Cin);
   ix641 : inv01 port map ( Y=>nx640, A=>A(16));
   ix173 : xnor2 port map ( Y=>nx172, A0=>A(17), A1=>nx643);
   ix644 : xnor2 port map ( Y=>nx643, A0=>B(17), A1=>Cin);
   ix648 : xnor2 port map ( Y=>nx647, A0=>B(18), A1=>Cin);
   ix650 : inv01 port map ( Y=>nx649, A=>A(18));
   ix193 : xnor2 port map ( Y=>nx192, A0=>A(19), A1=>nx652);
   ix653 : xnor2 port map ( Y=>nx652, A0=>B(19), A1=>Cin);
   ix657 : xnor2 port map ( Y=>nx656, A0=>B(20), A1=>Cin);
   ix659 : inv01 port map ( Y=>nx658, A=>A(20));
   ix213 : xnor2 port map ( Y=>nx212, A0=>A(21), A1=>nx661);
   ix662 : xnor2 port map ( Y=>nx661, A0=>B(21), A1=>Cin);
   ix666 : xnor2 port map ( Y=>nx665, A0=>B(22), A1=>Cin);
   ix668 : inv01 port map ( Y=>nx667, A=>A(22));
   ix233 : xnor2 port map ( Y=>nx232, A0=>A(23), A1=>nx670);
   ix671 : xnor2 port map ( Y=>nx670, A0=>B(23), A1=>Cin);
   ix675 : xnor2 port map ( Y=>nx674, A0=>B(24), A1=>Cin);
   ix677 : inv01 port map ( Y=>nx676, A=>A(24));
   ix253 : xnor2 port map ( Y=>nx252, A0=>A(25), A1=>nx679);
   ix680 : xnor2 port map ( Y=>nx679, A0=>B(25), A1=>Cin);
   ix684 : xnor2 port map ( Y=>nx683, A0=>B(26), A1=>Cin);
   ix686 : inv01 port map ( Y=>nx685, A=>A(26));
   ix273 : xnor2 port map ( Y=>nx272, A0=>A(27), A1=>nx688);
   ix689 : xnor2 port map ( Y=>nx688, A0=>B(27), A1=>Cin);
   ix693 : xnor2 port map ( Y=>nx692, A0=>B(28), A1=>Cin);
   ix695 : inv01 port map ( Y=>nx694, A=>A(28));
   ix293 : xnor2 port map ( Y=>nx292, A0=>A(29), A1=>nx697);
   ix698 : xnor2 port map ( Y=>nx697, A0=>B(29), A1=>Cin);
   ix702 : xnor2 port map ( Y=>nx701, A0=>B(30), A1=>Cin);
   ix704 : inv01 port map ( Y=>nx703, A=>A(30));
   ix313 : xnor2 port map ( Y=>nx312, A0=>A(31), A1=>nx706);
   ix707 : xnor2 port map ( Y=>nx706, A0=>B(31), A1=>Cin);
   ix383 : xor2 port map ( Y=>Sum(0), A0=>A(0), A1=>B(0));
   ix381 : xor2 port map ( Y=>Sum(1), A0=>nx8, A1=>nx12);
   ix379 : xnor2 port map ( Y=>Sum(2), A0=>nx566, A1=>nx22);
   ix23 : xnor2 port map ( Y=>nx22, A0=>A(2), A1=>nx575);
   ix377 : xor2 port map ( Y=>Sum(3), A0=>nx28, A1=>nx32);
   ix375 : xnor2 port map ( Y=>Sum(4), A0=>nx562, A1=>nx42);
   ix43 : xnor2 port map ( Y=>nx42, A0=>A(4), A1=>nx584);
   ix373 : xor2 port map ( Y=>Sum(5), A0=>nx48, A1=>nx52);
   ix371 : xnor2 port map ( Y=>Sum(6), A0=>nx558, A1=>nx62);
   ix63 : xnor2 port map ( Y=>nx62, A0=>A(6), A1=>nx593);
   ix369 : xor2 port map ( Y=>Sum(7), A0=>nx68, A1=>nx72);
   ix367 : xnor2 port map ( Y=>Sum(8), A0=>nx554, A1=>nx82);
   ix83 : xnor2 port map ( Y=>nx82, A0=>A(8), A1=>nx602);
   ix365 : xor2 port map ( Y=>Sum(9), A0=>nx88, A1=>nx92);
   ix363 : xnor2 port map ( Y=>Sum(10), A0=>nx550, A1=>nx102);
   ix103 : xnor2 port map ( Y=>nx102, A0=>A(10), A1=>nx611);
   ix361 : xor2 port map ( Y=>Sum(11), A0=>nx108, A1=>nx112);
   ix359 : xnor2 port map ( Y=>Sum(12), A0=>nx546, A1=>nx122);
   ix123 : xnor2 port map ( Y=>nx122, A0=>A(12), A1=>nx620);
   ix357 : xor2 port map ( Y=>Sum(13), A0=>nx128, A1=>nx132);
   ix355 : xnor2 port map ( Y=>Sum(14), A0=>nx542, A1=>nx142);
   ix143 : xnor2 port map ( Y=>nx142, A0=>A(14), A1=>nx629);
   ix353 : xor2 port map ( Y=>Sum(15), A0=>nx148, A1=>nx152);
   ix351 : xnor2 port map ( Y=>Sum(16), A0=>nx538, A1=>nx162);
   ix163 : xnor2 port map ( Y=>nx162, A0=>A(16), A1=>nx638);
   ix349 : xor2 port map ( Y=>Sum(17), A0=>nx168, A1=>nx172);
   ix347 : xnor2 port map ( Y=>Sum(18), A0=>nx534, A1=>nx182);
   ix183 : xnor2 port map ( Y=>nx182, A0=>A(18), A1=>nx647);
   ix345 : xor2 port map ( Y=>Sum(19), A0=>nx188, A1=>nx192);
   ix343 : xnor2 port map ( Y=>Sum(20), A0=>nx530, A1=>nx202);
   ix203 : xnor2 port map ( Y=>nx202, A0=>A(20), A1=>nx656);
   ix341 : xor2 port map ( Y=>Sum(21), A0=>nx208, A1=>nx212);
   ix339 : xnor2 port map ( Y=>Sum(22), A0=>nx526, A1=>nx222);
   ix223 : xnor2 port map ( Y=>nx222, A0=>A(22), A1=>nx665);
   ix337 : xor2 port map ( Y=>Sum(23), A0=>nx228, A1=>nx232);
   ix335 : xnor2 port map ( Y=>Sum(24), A0=>nx522, A1=>nx242);
   ix243 : xnor2 port map ( Y=>nx242, A0=>A(24), A1=>nx674);
   ix333 : xor2 port map ( Y=>Sum(25), A0=>nx248, A1=>nx252);
   ix331 : xnor2 port map ( Y=>Sum(26), A0=>nx518, A1=>nx262);
   ix263 : xnor2 port map ( Y=>nx262, A0=>A(26), A1=>nx683);
   ix329 : xor2 port map ( Y=>Sum(27), A0=>nx268, A1=>nx272);
   ix327 : xnor2 port map ( Y=>Sum(28), A0=>nx514, A1=>nx282);
   ix283 : xnor2 port map ( Y=>nx282, A0=>A(28), A1=>nx692);
   ix325 : xor2 port map ( Y=>Sum(29), A0=>nx288, A1=>nx292);
   ix323 : xnor2 port map ( Y=>Sum(30), A0=>nx510, A1=>nx302);
   ix303 : xnor2 port map ( Y=>nx302, A0=>A(30), A1=>nx701);
   ix315 : xor2 port map ( Y=>Sum(31), A0=>nx308, A1=>nx312);
   ix311 : inv01 port map ( Y=>nx310, A=>nx706);
   ix700 : inv01 port map ( Y=>nx699, A=>nx302);
   ix291 : inv01 port map ( Y=>nx290, A=>nx697);
   ix691 : inv01 port map ( Y=>nx690, A=>nx282);
   ix271 : inv01 port map ( Y=>nx270, A=>nx688);
   ix682 : inv01 port map ( Y=>nx681, A=>nx262);
   ix251 : inv01 port map ( Y=>nx250, A=>nx679);
   ix673 : inv01 port map ( Y=>nx672, A=>nx242);
   ix231 : inv01 port map ( Y=>nx230, A=>nx670);
   ix664 : inv01 port map ( Y=>nx663, A=>nx222);
   ix211 : inv01 port map ( Y=>nx210, A=>nx661);
   ix655 : inv01 port map ( Y=>nx654, A=>nx202);
   ix191 : inv01 port map ( Y=>nx190, A=>nx652);
   ix646 : inv01 port map ( Y=>nx645, A=>nx182);
   ix171 : inv01 port map ( Y=>nx170, A=>nx643);
   ix637 : inv01 port map ( Y=>nx636, A=>nx162);
   ix151 : inv01 port map ( Y=>nx150, A=>nx634);
   ix628 : inv01 port map ( Y=>nx627, A=>nx142);
   ix131 : inv01 port map ( Y=>nx130, A=>nx625);
   ix619 : inv01 port map ( Y=>nx618, A=>nx122);
   ix111 : inv01 port map ( Y=>nx110, A=>nx616);
   ix610 : inv01 port map ( Y=>nx609, A=>nx102);
   ix91 : inv01 port map ( Y=>nx90, A=>nx607);
   ix601 : inv01 port map ( Y=>nx600, A=>nx82);
   ix71 : inv01 port map ( Y=>nx70, A=>nx598);
   ix592 : inv01 port map ( Y=>nx591, A=>nx62);
   ix51 : inv01 port map ( Y=>nx50, A=>nx589);
   ix583 : inv01 port map ( Y=>nx582, A=>nx42);
   ix31 : inv01 port map ( Y=>nx30, A=>nx580);
   ix574 : inv01 port map ( Y=>nx573, A=>nx22);
   ix11 : inv01 port map ( Y=>nx10, A=>nx571);
end structural ;

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity RegisterN_32 is
   port (
      clk : IN std_logic ;
      reset : IN std_logic ;
      enable : IN std_logic ;
      input : IN std_logic_vector (31 DOWNTO 0) ;
      output : OUT std_logic_vector (31 DOWNTO 0)) ;
end RegisterN_32 ;

architecture Behavioral of RegisterN_32 is
   signal output_31_EXMPLR, output_30_EXMPLR, output_29_EXMPLR, 
      output_28_EXMPLR, output_27_EXMPLR, output_26_EXMPLR, output_25_EXMPLR, 
      output_24_EXMPLR, output_23_EXMPLR, output_22_EXMPLR, output_21_EXMPLR, 
      output_20_EXMPLR, output_19_EXMPLR, output_18_EXMPLR, output_17_EXMPLR, 
      output_16_EXMPLR, output_15_EXMPLR, output_14_EXMPLR, output_13_EXMPLR, 
      output_12_EXMPLR, output_11_EXMPLR, output_10_EXMPLR, output_9_EXMPLR, 
      output_8_EXMPLR, output_7_EXMPLR, output_6_EXMPLR, output_5_EXMPLR, 
      output_4_EXMPLR, output_3_EXMPLR, output_2_EXMPLR, output_1_EXMPLR, 
      output_0_EXMPLR, NOT_reset, nx422, nx432, nx442, nx452, nx462, nx472, 
      nx482, nx492, nx502, nx512, nx522, nx532, nx542, nx552, nx562, nx572, 
      nx582, nx592, nx602, nx612, nx622, nx632, nx642, nx652, nx662, nx672, 
      nx682, nx692, nx702, nx712, nx722, nx732, nx845, nx847: std_logic ;

begin
   output(31) <= output_31_EXMPLR ;
   output(30) <= output_30_EXMPLR ;
   output(29) <= output_29_EXMPLR ;
   output(28) <= output_28_EXMPLR ;
   output(27) <= output_27_EXMPLR ;
   output(26) <= output_26_EXMPLR ;
   output(25) <= output_25_EXMPLR ;
   output(24) <= output_24_EXMPLR ;
   output(23) <= output_23_EXMPLR ;
   output(22) <= output_22_EXMPLR ;
   output(21) <= output_21_EXMPLR ;
   output(20) <= output_20_EXMPLR ;
   output(19) <= output_19_EXMPLR ;
   output(18) <= output_18_EXMPLR ;
   output(17) <= output_17_EXMPLR ;
   output(16) <= output_16_EXMPLR ;
   output(15) <= output_15_EXMPLR ;
   output(14) <= output_14_EXMPLR ;
   output(13) <= output_13_EXMPLR ;
   output(12) <= output_12_EXMPLR ;
   output(11) <= output_11_EXMPLR ;
   output(10) <= output_10_EXMPLR ;
   output(9) <= output_9_EXMPLR ;
   output(8) <= output_8_EXMPLR ;
   output(7) <= output_7_EXMPLR ;
   output(6) <= output_6_EXMPLR ;
   output(5) <= output_5_EXMPLR ;
   output(4) <= output_4_EXMPLR ;
   output(3) <= output_3_EXMPLR ;
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   reg_output_0 : dffr port map ( Q=>output_0_EXMPLR, QB=>OPEN, D=>nx422, 
      CLK=>clk, R=>nx845);
   ix423 : mux21 port map ( Y=>nx422, A0=>output_0_EXMPLR, A1=>input(0), S0
      =>enable);
   ix745 : inv01 port map ( Y=>NOT_reset, A=>reset);
   reg_output_1 : dffr port map ( Q=>output_1_EXMPLR, QB=>OPEN, D=>nx432, 
      CLK=>clk, R=>nx845);
   ix433 : mux21 port map ( Y=>nx432, A0=>output_1_EXMPLR, A1=>input(1), S0
      =>enable);
   reg_output_2 : dffr port map ( Q=>output_2_EXMPLR, QB=>OPEN, D=>nx442, 
      CLK=>clk, R=>nx845);
   ix443 : mux21 port map ( Y=>nx442, A0=>output_2_EXMPLR, A1=>input(2), S0
      =>enable);
   reg_output_3 : dffr port map ( Q=>output_3_EXMPLR, QB=>OPEN, D=>nx452, 
      CLK=>clk, R=>nx845);
   ix453 : mux21 port map ( Y=>nx452, A0=>output_3_EXMPLR, A1=>input(3), S0
      =>enable);
   reg_output_4 : dffr port map ( Q=>output_4_EXMPLR, QB=>OPEN, D=>nx462, 
      CLK=>clk, R=>nx845);
   ix463 : mux21 port map ( Y=>nx462, A0=>output_4_EXMPLR, A1=>input(4), S0
      =>enable);
   reg_output_5 : dffr port map ( Q=>output_5_EXMPLR, QB=>OPEN, D=>nx472, 
      CLK=>clk, R=>nx845);
   ix473 : mux21 port map ( Y=>nx472, A0=>output_5_EXMPLR, A1=>input(5), S0
      =>enable);
   reg_output_6 : dffr port map ( Q=>output_6_EXMPLR, QB=>OPEN, D=>nx482, 
      CLK=>clk, R=>nx845);
   ix483 : mux21 port map ( Y=>nx482, A0=>output_6_EXMPLR, A1=>input(6), S0
      =>enable);
   reg_output_7 : dffr port map ( Q=>output_7_EXMPLR, QB=>OPEN, D=>nx492, 
      CLK=>clk, R=>nx845);
   ix493 : mux21 port map ( Y=>nx492, A0=>output_7_EXMPLR, A1=>input(7), S0
      =>enable);
   reg_output_8 : dffr port map ( Q=>output_8_EXMPLR, QB=>OPEN, D=>nx502, 
      CLK=>clk, R=>nx845);
   ix503 : mux21 port map ( Y=>nx502, A0=>output_8_EXMPLR, A1=>input(8), S0
      =>enable);
   reg_output_9 : dffr port map ( Q=>output_9_EXMPLR, QB=>OPEN, D=>nx512, 
      CLK=>clk, R=>nx845);
   ix513 : mux21 port map ( Y=>nx512, A0=>output_9_EXMPLR, A1=>input(9), S0
      =>enable);
   reg_output_10 : dffr port map ( Q=>output_10_EXMPLR, QB=>OPEN, D=>nx522, 
      CLK=>clk, R=>nx845);
   ix523 : mux21 port map ( Y=>nx522, A0=>output_10_EXMPLR, A1=>input(10), 
      S0=>enable);
   reg_output_11 : dffr port map ( Q=>output_11_EXMPLR, QB=>OPEN, D=>nx532, 
      CLK=>clk, R=>nx845);
   ix533 : mux21 port map ( Y=>nx532, A0=>output_11_EXMPLR, A1=>input(11), 
      S0=>enable);
   reg_output_12 : dffr port map ( Q=>output_12_EXMPLR, QB=>OPEN, D=>nx542, 
      CLK=>clk, R=>nx845);
   ix543 : mux21 port map ( Y=>nx542, A0=>output_12_EXMPLR, A1=>input(12), 
      S0=>enable);
   reg_output_13 : dffr port map ( Q=>output_13_EXMPLR, QB=>OPEN, D=>nx552, 
      CLK=>clk, R=>nx845);
   ix553 : mux21 port map ( Y=>nx552, A0=>output_13_EXMPLR, A1=>input(13), 
      S0=>enable);
   reg_output_14 : dffr port map ( Q=>output_14_EXMPLR, QB=>OPEN, D=>nx562, 
      CLK=>clk, R=>nx845);
   ix563 : mux21 port map ( Y=>nx562, A0=>output_14_EXMPLR, A1=>input(14), 
      S0=>enable);
   reg_output_15 : dffr port map ( Q=>output_15_EXMPLR, QB=>OPEN, D=>nx572, 
      CLK=>clk, R=>nx847);
   ix573 : mux21 port map ( Y=>nx572, A0=>output_15_EXMPLR, A1=>input(15), 
      S0=>enable);
   reg_output_16 : dffr port map ( Q=>output_16_EXMPLR, QB=>OPEN, D=>nx582, 
      CLK=>clk, R=>nx847);
   ix583 : mux21 port map ( Y=>nx582, A0=>output_16_EXMPLR, A1=>input(16), 
      S0=>enable);
   reg_output_17 : dffr port map ( Q=>output_17_EXMPLR, QB=>OPEN, D=>nx592, 
      CLK=>clk, R=>nx847);
   ix593 : mux21 port map ( Y=>nx592, A0=>output_17_EXMPLR, A1=>input(17), 
      S0=>enable);
   reg_output_18 : dffr port map ( Q=>output_18_EXMPLR, QB=>OPEN, D=>nx602, 
      CLK=>clk, R=>nx847);
   ix603 : mux21 port map ( Y=>nx602, A0=>output_18_EXMPLR, A1=>input(18), 
      S0=>enable);
   reg_output_19 : dffr port map ( Q=>output_19_EXMPLR, QB=>OPEN, D=>nx612, 
      CLK=>clk, R=>nx847);
   ix613 : mux21 port map ( Y=>nx612, A0=>output_19_EXMPLR, A1=>input(19), 
      S0=>enable);
   reg_output_20 : dffr port map ( Q=>output_20_EXMPLR, QB=>OPEN, D=>nx622, 
      CLK=>clk, R=>nx847);
   ix623 : mux21 port map ( Y=>nx622, A0=>output_20_EXMPLR, A1=>input(20), 
      S0=>enable);
   reg_output_21 : dffr port map ( Q=>output_21_EXMPLR, QB=>OPEN, D=>nx632, 
      CLK=>clk, R=>nx847);
   ix633 : mux21 port map ( Y=>nx632, A0=>output_21_EXMPLR, A1=>input(21), 
      S0=>enable);
   reg_output_22 : dffr port map ( Q=>output_22_EXMPLR, QB=>OPEN, D=>nx642, 
      CLK=>clk, R=>nx847);
   ix643 : mux21 port map ( Y=>nx642, A0=>output_22_EXMPLR, A1=>input(22), 
      S0=>enable);
   reg_output_23 : dffr port map ( Q=>output_23_EXMPLR, QB=>OPEN, D=>nx652, 
      CLK=>clk, R=>nx847);
   ix653 : mux21 port map ( Y=>nx652, A0=>output_23_EXMPLR, A1=>input(23), 
      S0=>enable);
   reg_output_24 : dffr port map ( Q=>output_24_EXMPLR, QB=>OPEN, D=>nx662, 
      CLK=>clk, R=>nx847);
   ix663 : mux21 port map ( Y=>nx662, A0=>output_24_EXMPLR, A1=>input(24), 
      S0=>enable);
   reg_output_25 : dffr port map ( Q=>output_25_EXMPLR, QB=>OPEN, D=>nx672, 
      CLK=>clk, R=>nx847);
   ix673 : mux21 port map ( Y=>nx672, A0=>output_25_EXMPLR, A1=>input(25), 
      S0=>enable);
   reg_output_26 : dffr port map ( Q=>output_26_EXMPLR, QB=>OPEN, D=>nx682, 
      CLK=>clk, R=>nx847);
   ix683 : mux21 port map ( Y=>nx682, A0=>output_26_EXMPLR, A1=>input(26), 
      S0=>enable);
   reg_output_27 : dffr port map ( Q=>output_27_EXMPLR, QB=>OPEN, D=>nx692, 
      CLK=>clk, R=>nx847);
   ix693 : mux21 port map ( Y=>nx692, A0=>output_27_EXMPLR, A1=>input(27), 
      S0=>enable);
   reg_output_28 : dffr port map ( Q=>output_28_EXMPLR, QB=>OPEN, D=>nx702, 
      CLK=>clk, R=>nx847);
   ix703 : mux21 port map ( Y=>nx702, A0=>output_28_EXMPLR, A1=>input(28), 
      S0=>enable);
   reg_output_29 : dffr port map ( Q=>output_29_EXMPLR, QB=>OPEN, D=>nx712, 
      CLK=>clk, R=>nx847);
   ix713 : mux21 port map ( Y=>nx712, A0=>output_29_EXMPLR, A1=>input(29), 
      S0=>enable);
   reg_output_30 : dffr port map ( Q=>output_30_EXMPLR, QB=>OPEN, D=>nx722, 
      CLK=>clk, R=>NOT_reset);
   ix723 : mux21 port map ( Y=>nx722, A0=>output_30_EXMPLR, A1=>input(30), 
      S0=>enable);
   reg_output_31 : dffr port map ( Q=>output_31_EXMPLR, QB=>OPEN, D=>nx732, 
      CLK=>clk, R=>NOT_reset);
   ix733 : mux21 port map ( Y=>nx732, A0=>output_31_EXMPLR, A1=>input(31), 
      S0=>enable);
   ix844 : inv01 port map ( Y=>nx845, A=>reset);
   ix846 : inv01 port map ( Y=>nx847, A=>reset);
end Behavioral ;

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity LFSR is
   port (
      clk : IN std_logic ;
      rst : IN std_logic ;
      enable : IN std_logic ;
      bit_pattern : OUT std_logic_vector (31 DOWNTO 0)) ;
end LFSR ;

architecture Behavioral of LFSR is
   signal bit_pattern_31_EXMPLR, bit_pattern_30_EXMPLR, 
      bit_pattern_29_EXMPLR, bit_pattern_28_EXMPLR, bit_pattern_27_EXMPLR, 
      bit_pattern_26_EXMPLR, bit_pattern_25_EXMPLR, bit_pattern_24_EXMPLR, 
      bit_pattern_23_EXMPLR, bit_pattern_22_EXMPLR, bit_pattern_21_EXMPLR, 
      bit_pattern_20_EXMPLR, bit_pattern_19_EXMPLR, bit_pattern_18_EXMPLR, 
      bit_pattern_17_EXMPLR, bit_pattern_16_EXMPLR, bit_pattern_15_EXMPLR, 
      bit_pattern_14_EXMPLR, bit_pattern_13_EXMPLR, bit_pattern_12_EXMPLR, 
      bit_pattern_11_EXMPLR, bit_pattern_10_EXMPLR, bit_pattern_9_EXMPLR, 
      bit_pattern_8_EXMPLR, bit_pattern_7_EXMPLR, bit_pattern_6_EXMPLR, 
      bit_pattern_5_EXMPLR, bit_pattern_4_EXMPLR, bit_pattern_3_EXMPLR, 
      bit_pattern_2_EXMPLR, bit_pattern_1_EXMPLR, bit_pattern_0_EXMPLR, 
      zeroth_in, nx38, nx72, nx82, nx740, nx750, nx760, nx770, nx780, nx790, 
      nx800, nx810, nx820, nx830, nx840, nx850, nx860, nx870, nx880, nx890, 
      nx900, nx910, nx920, nx930, nx940, nx950, nx960, nx970, nx980, nx990, 
      nx1000, nx1010, nx1020, nx1030, nx1040, nx1050, nx1060, nx1139, nx1144, 
      nx1183, nx1185, nx1187, nx1189: std_logic ;

begin
   bit_pattern(31) <= bit_pattern_31_EXMPLR ;
   bit_pattern(30) <= bit_pattern_30_EXMPLR ;
   bit_pattern(29) <= bit_pattern_29_EXMPLR ;
   bit_pattern(28) <= bit_pattern_28_EXMPLR ;
   bit_pattern(27) <= bit_pattern_27_EXMPLR ;
   bit_pattern(26) <= bit_pattern_26_EXMPLR ;
   bit_pattern(25) <= bit_pattern_25_EXMPLR ;
   bit_pattern(24) <= bit_pattern_24_EXMPLR ;
   bit_pattern(23) <= bit_pattern_23_EXMPLR ;
   bit_pattern(22) <= bit_pattern_22_EXMPLR ;
   bit_pattern(21) <= bit_pattern_21_EXMPLR ;
   bit_pattern(20) <= bit_pattern_20_EXMPLR ;
   bit_pattern(19) <= bit_pattern_19_EXMPLR ;
   bit_pattern(18) <= bit_pattern_18_EXMPLR ;
   bit_pattern(17) <= bit_pattern_17_EXMPLR ;
   bit_pattern(16) <= bit_pattern_16_EXMPLR ;
   bit_pattern(15) <= bit_pattern_15_EXMPLR ;
   bit_pattern(14) <= bit_pattern_14_EXMPLR ;
   bit_pattern(13) <= bit_pattern_13_EXMPLR ;
   bit_pattern(12) <= bit_pattern_12_EXMPLR ;
   bit_pattern(11) <= bit_pattern_11_EXMPLR ;
   bit_pattern(10) <= bit_pattern_10_EXMPLR ;
   bit_pattern(9) <= bit_pattern_9_EXMPLR ;
   bit_pattern(8) <= bit_pattern_8_EXMPLR ;
   bit_pattern(7) <= bit_pattern_7_EXMPLR ;
   bit_pattern(6) <= bit_pattern_6_EXMPLR ;
   bit_pattern(5) <= bit_pattern_5_EXMPLR ;
   bit_pattern(4) <= bit_pattern_4_EXMPLR ;
   bit_pattern(3) <= bit_pattern_3_EXMPLR ;
   bit_pattern(2) <= bit_pattern_2_EXMPLR ;
   bit_pattern(1) <= bit_pattern_1_EXMPLR ;
   bit_pattern(0) <= bit_pattern_0_EXMPLR ;
   reg_LFSR_REG_0 : dff port map ( Q=>bit_pattern_0_EXMPLR, QB=>OPEN, D=>
      nx740, CLK=>clk);
   ix741 : ao221 port map ( Y=>nx740, A0=>bit_pattern_1_EXMPLR, A1=>enable, 
      B0=>bit_pattern_0_EXMPLR, B1=>nx1189, C0=>nx1144);
   reg_LFSR_REG_1 : dff port map ( Q=>bit_pattern_1_EXMPLR, QB=>OPEN, D=>
      nx1060, CLK=>clk);
   ix1061 : ao32 port map ( Y=>nx1060, A0=>rst, A1=>bit_pattern_2_EXMPLR, A2
      =>enable, B0=>bit_pattern_1_EXMPLR, B1=>nx1189);
   reg_LFSR_REG_2 : dff port map ( Q=>bit_pattern_2_EXMPLR, QB=>OPEN, D=>
      nx1050, CLK=>clk);
   ix1051 : ao32 port map ( Y=>nx1050, A0=>rst, A1=>bit_pattern_3_EXMPLR, A2
      =>enable, B0=>bit_pattern_2_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_3 : dff port map ( Q=>bit_pattern_3_EXMPLR, QB=>OPEN, D=>
      nx1040, CLK=>clk);
   ix1041 : ao32 port map ( Y=>nx1040, A0=>rst, A1=>bit_pattern_4_EXMPLR, A2
      =>enable, B0=>bit_pattern_3_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_4 : dff port map ( Q=>bit_pattern_4_EXMPLR, QB=>OPEN, D=>
      nx1030, CLK=>clk);
   ix1031 : ao32 port map ( Y=>nx1030, A0=>rst, A1=>bit_pattern_5_EXMPLR, A2
      =>enable, B0=>bit_pattern_4_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_5 : dff port map ( Q=>bit_pattern_5_EXMPLR, QB=>OPEN, D=>
      nx1020, CLK=>clk);
   ix1021 : ao32 port map ( Y=>nx1020, A0=>rst, A1=>bit_pattern_6_EXMPLR, A2
      =>enable, B0=>bit_pattern_5_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_6 : dff port map ( Q=>bit_pattern_6_EXMPLR, QB=>OPEN, D=>
      nx1010, CLK=>clk);
   ix1011 : ao32 port map ( Y=>nx1010, A0=>rst, A1=>bit_pattern_7_EXMPLR, A2
      =>enable, B0=>bit_pattern_6_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_7 : dff port map ( Q=>bit_pattern_7_EXMPLR, QB=>OPEN, D=>
      nx1000, CLK=>clk);
   ix1001 : ao32 port map ( Y=>nx1000, A0=>rst, A1=>bit_pattern_8_EXMPLR, A2
      =>enable, B0=>bit_pattern_7_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_8 : dff port map ( Q=>bit_pattern_8_EXMPLR, QB=>OPEN, D=>
      nx990, CLK=>clk);
   ix991 : ao32 port map ( Y=>nx990, A0=>rst, A1=>bit_pattern_9_EXMPLR, A2=>
      enable, B0=>bit_pattern_8_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_9 : dff port map ( Q=>bit_pattern_9_EXMPLR, QB=>OPEN, D=>
      nx980, CLK=>clk);
   ix981 : ao32 port map ( Y=>nx980, A0=>rst, A1=>bit_pattern_10_EXMPLR, A2
      =>enable, B0=>bit_pattern_9_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_10 : dff port map ( Q=>bit_pattern_10_EXMPLR, QB=>OPEN, D=>
      nx970, CLK=>clk);
   ix971 : ao32 port map ( Y=>nx970, A0=>rst, A1=>bit_pattern_11_EXMPLR, A2
      =>enable, B0=>bit_pattern_10_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_11 : dff port map ( Q=>bit_pattern_11_EXMPLR, QB=>OPEN, D=>
      nx960, CLK=>clk);
   ix961 : ao32 port map ( Y=>nx960, A0=>rst, A1=>bit_pattern_12_EXMPLR, A2
      =>enable, B0=>bit_pattern_11_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_12 : dff port map ( Q=>bit_pattern_12_EXMPLR, QB=>OPEN, D=>
      nx950, CLK=>clk);
   ix951 : ao32 port map ( Y=>nx950, A0=>rst, A1=>bit_pattern_13_EXMPLR, A2
      =>enable, B0=>bit_pattern_12_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_13 : dff port map ( Q=>bit_pattern_13_EXMPLR, QB=>OPEN, D=>
      nx940, CLK=>clk);
   ix941 : ao32 port map ( Y=>nx940, A0=>rst, A1=>bit_pattern_14_EXMPLR, A2
      =>enable, B0=>bit_pattern_13_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_14 : dff port map ( Q=>bit_pattern_14_EXMPLR, QB=>OPEN, D=>
      nx930, CLK=>clk);
   ix931 : ao32 port map ( Y=>nx930, A0=>rst, A1=>bit_pattern_15_EXMPLR, A2
      =>enable, B0=>bit_pattern_14_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_15 : dff port map ( Q=>bit_pattern_15_EXMPLR, QB=>OPEN, D=>
      nx920, CLK=>clk);
   ix921 : ao32 port map ( Y=>nx920, A0=>rst, A1=>bit_pattern_16_EXMPLR, A2
      =>enable, B0=>bit_pattern_15_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_16 : dff port map ( Q=>bit_pattern_16_EXMPLR, QB=>OPEN, D=>
      nx910, CLK=>clk);
   ix911 : ao32 port map ( Y=>nx910, A0=>rst, A1=>bit_pattern_17_EXMPLR, A2
      =>enable, B0=>bit_pattern_16_EXMPLR, B1=>nx1187);
   reg_LFSR_REG_17 : dff port map ( Q=>bit_pattern_17_EXMPLR, QB=>OPEN, D=>
      nx900, CLK=>clk);
   ix901 : ao32 port map ( Y=>nx900, A0=>rst, A1=>bit_pattern_18_EXMPLR, A2
      =>enable, B0=>bit_pattern_17_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_18 : dff port map ( Q=>bit_pattern_18_EXMPLR, QB=>OPEN, D=>
      nx890, CLK=>clk);
   ix891 : ao32 port map ( Y=>nx890, A0=>rst, A1=>bit_pattern_19_EXMPLR, A2
      =>enable, B0=>bit_pattern_18_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_19 : dff port map ( Q=>bit_pattern_19_EXMPLR, QB=>OPEN, D=>
      nx880, CLK=>clk);
   ix881 : ao32 port map ( Y=>nx880, A0=>rst, A1=>bit_pattern_20_EXMPLR, A2
      =>enable, B0=>bit_pattern_19_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_20 : dff port map ( Q=>bit_pattern_20_EXMPLR, QB=>OPEN, D=>
      nx870, CLK=>clk);
   ix871 : ao32 port map ( Y=>nx870, A0=>rst, A1=>bit_pattern_21_EXMPLR, A2
      =>enable, B0=>bit_pattern_20_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_21 : dff port map ( Q=>bit_pattern_21_EXMPLR, QB=>OPEN, D=>
      nx860, CLK=>clk);
   ix861 : ao32 port map ( Y=>nx860, A0=>rst, A1=>bit_pattern_22_EXMPLR, A2
      =>enable, B0=>bit_pattern_21_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_22 : dff port map ( Q=>bit_pattern_22_EXMPLR, QB=>OPEN, D=>
      nx850, CLK=>clk);
   ix851 : ao32 port map ( Y=>nx850, A0=>rst, A1=>bit_pattern_23_EXMPLR, A2
      =>enable, B0=>bit_pattern_22_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_23 : dff port map ( Q=>bit_pattern_23_EXMPLR, QB=>OPEN, D=>
      nx840, CLK=>clk);
   ix841 : ao32 port map ( Y=>nx840, A0=>rst, A1=>bit_pattern_24_EXMPLR, A2
      =>enable, B0=>bit_pattern_23_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_24 : dff port map ( Q=>bit_pattern_24_EXMPLR, QB=>OPEN, D=>
      nx830, CLK=>clk);
   ix831 : ao32 port map ( Y=>nx830, A0=>rst, A1=>nx82, A2=>enable, B0=>
      bit_pattern_24_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_25 : dff port map ( Q=>bit_pattern_25_EXMPLR, QB=>OPEN, D=>
      nx820, CLK=>clk);
   ix821 : ao32 port map ( Y=>nx820, A0=>rst, A1=>nx72, A2=>enable, B0=>
      bit_pattern_25_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_26 : dff port map ( Q=>bit_pattern_26_EXMPLR, QB=>OPEN, D=>
      nx810, CLK=>clk);
   ix811 : ao32 port map ( Y=>nx810, A0=>rst, A1=>bit_pattern_27_EXMPLR, A2
      =>enable, B0=>bit_pattern_26_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_27 : dff port map ( Q=>bit_pattern_27_EXMPLR, QB=>OPEN, D=>
      nx800, CLK=>clk);
   ix801 : ao32 port map ( Y=>nx800, A0=>rst, A1=>bit_pattern_28_EXMPLR, A2
      =>enable, B0=>bit_pattern_27_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_28 : dff port map ( Q=>bit_pattern_28_EXMPLR, QB=>OPEN, D=>
      nx790, CLK=>clk);
   ix791 : ao32 port map ( Y=>nx790, A0=>rst, A1=>bit_pattern_29_EXMPLR, A2
      =>enable, B0=>bit_pattern_28_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_29 : dff port map ( Q=>bit_pattern_29_EXMPLR, QB=>OPEN, D=>
      nx780, CLK=>clk);
   ix781 : ao32 port map ( Y=>nx780, A0=>rst, A1=>nx38, A2=>enable, B0=>
      bit_pattern_29_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_30 : dff port map ( Q=>bit_pattern_30_EXMPLR, QB=>OPEN, D=>
      nx770, CLK=>clk);
   ix771 : ao32 port map ( Y=>nx770, A0=>rst, A1=>bit_pattern_31_EXMPLR, A2
      =>enable, B0=>bit_pattern_30_EXMPLR, B1=>nx1185);
   reg_LFSR_REG_31 : dff port map ( Q=>bit_pattern_31_EXMPLR, QB=>OPEN, D=>
      nx760, CLK=>clk);
   ix761 : ao32 port map ( Y=>nx760, A0=>rst, A1=>zeroth_in, A2=>enable, B0
      =>bit_pattern_31_EXMPLR, B1=>nx1185);
   reg_zeroth_in : dff port map ( Q=>zeroth_in, QB=>OPEN, D=>nx750, CLK=>clk
   );
   ix751 : mux21 port map ( Y=>nx750, A0=>bit_pattern_0_EXMPLR, A1=>
      zeroth_in, S0=>nx1139);
   ix1140 : nand02 port map ( Y=>nx1139, A0=>enable, A1=>rst);
   ix1145 : inv01 port map ( Y=>nx1144, A=>rst);
   ix1184 : inv01 port map ( Y=>nx1185, A=>nx1183);
   ix1186 : inv01 port map ( Y=>nx1187, A=>nx1183);
   ix1188 : inv01 port map ( Y=>nx1189, A=>nx1183);
   ix83 : xor2 port map ( Y=>nx82, A0=>bit_pattern_25_EXMPLR, A1=>zeroth_in
   );
   ix73 : xor2 port map ( Y=>nx72, A0=>bit_pattern_26_EXMPLR, A1=>zeroth_in
   );
   ix39 : xor2 port map ( Y=>nx38, A0=>bit_pattern_30_EXMPLR, A1=>zeroth_in
   );
   ix1143 : or02 port map ( Y=>nx1183, A0=>nx1144, A1=>enable);
end Behavioral ;

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity MISR is
   port (
      clk : IN std_logic ;
      rst : IN std_logic ;
      enable : IN std_logic ;
      mult_result : IN std_logic_vector (31 DOWNTO 0) ;
      signature : OUT std_logic_vector (31 DOWNTO 0)) ;
end MISR ;

architecture Behavioral of MISR is
   signal signature_31_EXMPLR, signature_30_EXMPLR, signature_29_EXMPLR, 
      signature_28_EXMPLR, signature_27_EXMPLR, signature_26_EXMPLR, 
      signature_25_EXMPLR, signature_24_EXMPLR, signature_23_EXMPLR, 
      signature_22_EXMPLR, signature_21_EXMPLR, signature_20_EXMPLR, 
      signature_19_EXMPLR, signature_18_EXMPLR, signature_17_EXMPLR, 
      signature_16_EXMPLR, signature_15_EXMPLR, signature_14_EXMPLR, 
      signature_13_EXMPLR, signature_12_EXMPLR, signature_11_EXMPLR, 
      signature_10_EXMPLR, signature_9_EXMPLR, signature_8_EXMPLR, 
      signature_7_EXMPLR, signature_6_EXMPLR, signature_5_EXMPLR, 
      signature_4_EXMPLR, signature_3_EXMPLR, signature_2_EXMPLR, 
      signature_1_EXMPLR, signature_0_EXMPLR, zeroth_in, nx12, nx22, nx34, 
      nx44, nx54, nx64, nx76, nx88, nx98, nx108, nx118, nx128, nx138, nx148, 
      nx158, nx168, nx178, nx188, nx198, nx208, nx218, nx228, nx238, nx248, 
      nx258, nx268, nx278, nx288, nx298, nx308, nx318, nx328, nx836, nx846, 
      nx856, nx866, nx876, nx886, nx896, nx906, nx916, nx926, nx936, nx946, 
      nx956, nx966, nx976, nx986, nx996, nx1006, nx1016, nx1026, nx1036, 
      nx1046, nx1056, nx1066, nx1076, nx1086, nx1096, nx1106, nx1116, nx1126, 
      nx1136, nx1146, nx1156, nx1168, nx1170, nx1245, nx1250, nx1264, nx1272, 
      nx1276, nx1315, nx1317, nx1323, nx1325, nx1327, nx1329: std_logic ;

begin
   signature(31) <= signature_31_EXMPLR ;
   signature(30) <= signature_30_EXMPLR ;
   signature(29) <= signature_29_EXMPLR ;
   signature(28) <= signature_28_EXMPLR ;
   signature(27) <= signature_27_EXMPLR ;
   signature(26) <= signature_26_EXMPLR ;
   signature(25) <= signature_25_EXMPLR ;
   signature(24) <= signature_24_EXMPLR ;
   signature(23) <= signature_23_EXMPLR ;
   signature(22) <= signature_22_EXMPLR ;
   signature(21) <= signature_21_EXMPLR ;
   signature(20) <= signature_20_EXMPLR ;
   signature(19) <= signature_19_EXMPLR ;
   signature(18) <= signature_18_EXMPLR ;
   signature(17) <= signature_17_EXMPLR ;
   signature(16) <= signature_16_EXMPLR ;
   signature(15) <= signature_15_EXMPLR ;
   signature(14) <= signature_14_EXMPLR ;
   signature(13) <= signature_13_EXMPLR ;
   signature(12) <= signature_12_EXMPLR ;
   signature(11) <= signature_11_EXMPLR ;
   signature(10) <= signature_10_EXMPLR ;
   signature(9) <= signature_9_EXMPLR ;
   signature(8) <= signature_8_EXMPLR ;
   signature(7) <= signature_7_EXMPLR ;
   signature(6) <= signature_6_EXMPLR ;
   signature(5) <= signature_5_EXMPLR ;
   signature(4) <= signature_4_EXMPLR ;
   signature(3) <= signature_3_EXMPLR ;
   signature(2) <= signature_2_EXMPLR ;
   signature(1) <= signature_1_EXMPLR ;
   signature(0) <= signature_0_EXMPLR ;
   reg_MISR_REG_0 : dff port map ( Q=>signature_0_EXMPLR, QB=>OPEN, D=>
      nx1156, CLK=>clk);
   ix1157 : ao221 port map ( Y=>nx1156, A0=>signature_0_EXMPLR, A1=>nx1315, 
      B0=>nx328, B1=>nx1329, C0=>nx1170);
   ix1171 : inv01 port map ( Y=>nx1170, A=>rst);
   ix329 : xor2 port map ( Y=>nx328, A0=>mult_result(0), A1=>
      signature_1_EXMPLR);
   reg_MISR_REG_1 : dff port map ( Q=>signature_1_EXMPLR, QB=>OPEN, D=>
      nx1146, CLK=>clk);
   ix1147 : ao32 port map ( Y=>nx1146, A0=>rst, A1=>nx318, A2=>nx1329, B0=>
      signature_1_EXMPLR, B1=>nx1168);
   ix319 : xor2 port map ( Y=>nx318, A0=>mult_result(1), A1=>
      signature_2_EXMPLR);
   reg_MISR_REG_2 : dff port map ( Q=>signature_2_EXMPLR, QB=>OPEN, D=>
      nx1136, CLK=>clk);
   ix1137 : ao32 port map ( Y=>nx1136, A0=>rst, A1=>nx308, A2=>nx1329, B0=>
      signature_2_EXMPLR, B1=>nx1168);
   ix309 : xor2 port map ( Y=>nx308, A0=>mult_result(2), A1=>
      signature_3_EXMPLR);
   reg_MISR_REG_3 : dff port map ( Q=>signature_3_EXMPLR, QB=>OPEN, D=>
      nx1126, CLK=>clk);
   ix1127 : ao32 port map ( Y=>nx1126, A0=>rst, A1=>nx298, A2=>nx1327, B0=>
      signature_3_EXMPLR, B1=>nx1168);
   ix299 : xor2 port map ( Y=>nx298, A0=>mult_result(3), A1=>
      signature_4_EXMPLR);
   reg_MISR_REG_4 : dff port map ( Q=>signature_4_EXMPLR, QB=>OPEN, D=>
      nx1116, CLK=>clk);
   ix1117 : ao32 port map ( Y=>nx1116, A0=>rst, A1=>nx288, A2=>nx1327, B0=>
      signature_4_EXMPLR, B1=>nx1317);
   ix289 : xor2 port map ( Y=>nx288, A0=>mult_result(4), A1=>
      signature_5_EXMPLR);
   reg_MISR_REG_5 : dff port map ( Q=>signature_5_EXMPLR, QB=>OPEN, D=>
      nx1106, CLK=>clk);
   ix1107 : ao32 port map ( Y=>nx1106, A0=>rst, A1=>nx278, A2=>nx1327, B0=>
      signature_5_EXMPLR, B1=>nx1317);
   ix279 : xor2 port map ( Y=>nx278, A0=>mult_result(5), A1=>
      signature_6_EXMPLR);
   reg_MISR_REG_6 : dff port map ( Q=>signature_6_EXMPLR, QB=>OPEN, D=>
      nx1096, CLK=>clk);
   ix1097 : ao32 port map ( Y=>nx1096, A0=>rst, A1=>nx268, A2=>nx1327, B0=>
      signature_6_EXMPLR, B1=>nx1317);
   ix269 : xor2 port map ( Y=>nx268, A0=>mult_result(6), A1=>
      signature_7_EXMPLR);
   reg_MISR_REG_7 : dff port map ( Q=>signature_7_EXMPLR, QB=>OPEN, D=>
      nx1086, CLK=>clk);
   ix1087 : ao32 port map ( Y=>nx1086, A0=>rst, A1=>nx258, A2=>nx1327, B0=>
      signature_7_EXMPLR, B1=>nx1317);
   ix259 : xor2 port map ( Y=>nx258, A0=>mult_result(7), A1=>
      signature_8_EXMPLR);
   reg_MISR_REG_8 : dff port map ( Q=>signature_8_EXMPLR, QB=>OPEN, D=>
      nx1076, CLK=>clk);
   ix1077 : ao32 port map ( Y=>nx1076, A0=>rst, A1=>nx248, A2=>nx1327, B0=>
      signature_8_EXMPLR, B1=>nx1317);
   ix249 : xor2 port map ( Y=>nx248, A0=>mult_result(8), A1=>
      signature_9_EXMPLR);
   reg_MISR_REG_9 : dff port map ( Q=>signature_9_EXMPLR, QB=>OPEN, D=>
      nx1066, CLK=>clk);
   ix1067 : ao32 port map ( Y=>nx1066, A0=>rst, A1=>nx238, A2=>nx1327, B0=>
      signature_9_EXMPLR, B1=>nx1317);
   ix239 : xor2 port map ( Y=>nx238, A0=>mult_result(9), A1=>
      signature_10_EXMPLR);
   reg_MISR_REG_10 : dff port map ( Q=>signature_10_EXMPLR, QB=>OPEN, D=>
      nx1056, CLK=>clk);
   ix1057 : ao32 port map ( Y=>nx1056, A0=>rst, A1=>nx228, A2=>nx1327, B0=>
      signature_10_EXMPLR, B1=>nx1317);
   ix229 : xor2 port map ( Y=>nx228, A0=>mult_result(10), A1=>
      signature_11_EXMPLR);
   reg_MISR_REG_11 : dff port map ( Q=>signature_11_EXMPLR, QB=>OPEN, D=>
      nx1046, CLK=>clk);
   ix1047 : ao32 port map ( Y=>nx1046, A0=>rst, A1=>nx218, A2=>nx1327, B0=>
      signature_11_EXMPLR, B1=>nx1317);
   ix219 : xor2 port map ( Y=>nx218, A0=>mult_result(11), A1=>
      signature_12_EXMPLR);
   reg_MISR_REG_12 : dff port map ( Q=>signature_12_EXMPLR, QB=>OPEN, D=>
      nx1036, CLK=>clk);
   ix1037 : ao32 port map ( Y=>nx1036, A0=>rst, A1=>nx208, A2=>nx1327, B0=>
      signature_12_EXMPLR, B1=>nx1317);
   ix209 : xor2 port map ( Y=>nx208, A0=>mult_result(12), A1=>
      signature_13_EXMPLR);
   reg_MISR_REG_13 : dff port map ( Q=>signature_13_EXMPLR, QB=>OPEN, D=>
      nx1026, CLK=>clk);
   ix1027 : ao32 port map ( Y=>nx1026, A0=>rst, A1=>nx198, A2=>nx1327, B0=>
      signature_13_EXMPLR, B1=>nx1317);
   ix199 : xor2 port map ( Y=>nx198, A0=>mult_result(13), A1=>
      signature_14_EXMPLR);
   reg_MISR_REG_14 : dff port map ( Q=>signature_14_EXMPLR, QB=>OPEN, D=>
      nx1016, CLK=>clk);
   ix1017 : ao32 port map ( Y=>nx1016, A0=>rst, A1=>nx188, A2=>nx1327, B0=>
      signature_14_EXMPLR, B1=>nx1317);
   ix189 : xor2 port map ( Y=>nx188, A0=>mult_result(14), A1=>
      signature_15_EXMPLR);
   reg_MISR_REG_15 : dff port map ( Q=>signature_15_EXMPLR, QB=>OPEN, D=>
      nx1006, CLK=>clk);
   ix1007 : ao32 port map ( Y=>nx1006, A0=>rst, A1=>nx178, A2=>nx1327, B0=>
      signature_15_EXMPLR, B1=>nx1317);
   ix179 : xor2 port map ( Y=>nx178, A0=>mult_result(15), A1=>
      signature_16_EXMPLR);
   reg_MISR_REG_16 : dff port map ( Q=>signature_16_EXMPLR, QB=>OPEN, D=>
      nx996, CLK=>clk);
   ix997 : ao32 port map ( Y=>nx996, A0=>rst, A1=>nx168, A2=>nx1327, B0=>
      signature_16_EXMPLR, B1=>nx1317);
   ix169 : xor2 port map ( Y=>nx168, A0=>mult_result(16), A1=>
      signature_17_EXMPLR);
   reg_MISR_REG_17 : dff port map ( Q=>signature_17_EXMPLR, QB=>OPEN, D=>
      nx986, CLK=>clk);
   ix987 : ao32 port map ( Y=>nx986, A0=>rst, A1=>nx158, A2=>nx1327, B0=>
      signature_17_EXMPLR, B1=>nx1317);
   ix159 : xor2 port map ( Y=>nx158, A0=>mult_result(17), A1=>
      signature_18_EXMPLR);
   reg_MISR_REG_18 : dff port map ( Q=>signature_18_EXMPLR, QB=>OPEN, D=>
      nx976, CLK=>clk);
   ix977 : ao32 port map ( Y=>nx976, A0=>rst, A1=>nx148, A2=>nx1325, B0=>
      signature_18_EXMPLR, B1=>nx1317);
   ix149 : xor2 port map ( Y=>nx148, A0=>mult_result(18), A1=>
      signature_19_EXMPLR);
   reg_MISR_REG_19 : dff port map ( Q=>signature_19_EXMPLR, QB=>OPEN, D=>
      nx966, CLK=>clk);
   ix967 : ao32 port map ( Y=>nx966, A0=>rst, A1=>nx138, A2=>nx1325, B0=>
      signature_19_EXMPLR, B1=>nx1315);
   ix139 : xor2 port map ( Y=>nx138, A0=>mult_result(19), A1=>
      signature_20_EXMPLR);
   reg_MISR_REG_20 : dff port map ( Q=>signature_20_EXMPLR, QB=>OPEN, D=>
      nx956, CLK=>clk);
   ix957 : ao32 port map ( Y=>nx956, A0=>rst, A1=>nx128, A2=>nx1325, B0=>
      signature_20_EXMPLR, B1=>nx1315);
   ix129 : xor2 port map ( Y=>nx128, A0=>mult_result(20), A1=>
      signature_21_EXMPLR);
   reg_MISR_REG_21 : dff port map ( Q=>signature_21_EXMPLR, QB=>OPEN, D=>
      nx946, CLK=>clk);
   ix947 : ao32 port map ( Y=>nx946, A0=>rst, A1=>nx118, A2=>nx1325, B0=>
      signature_21_EXMPLR, B1=>nx1315);
   ix119 : xor2 port map ( Y=>nx118, A0=>mult_result(21), A1=>
      signature_22_EXMPLR);
   reg_MISR_REG_22 : dff port map ( Q=>signature_22_EXMPLR, QB=>OPEN, D=>
      nx936, CLK=>clk);
   ix937 : ao32 port map ( Y=>nx936, A0=>rst, A1=>nx108, A2=>nx1325, B0=>
      signature_22_EXMPLR, B1=>nx1315);
   ix109 : xor2 port map ( Y=>nx108, A0=>mult_result(22), A1=>
      signature_23_EXMPLR);
   reg_MISR_REG_23 : dff port map ( Q=>signature_23_EXMPLR, QB=>OPEN, D=>
      nx926, CLK=>clk);
   ix927 : ao32 port map ( Y=>nx926, A0=>rst, A1=>nx98, A2=>nx1325, B0=>
      signature_23_EXMPLR, B1=>nx1315);
   ix99 : xor2 port map ( Y=>nx98, A0=>mult_result(23), A1=>
      signature_24_EXMPLR);
   reg_MISR_REG_24 : dff port map ( Q=>signature_24_EXMPLR, QB=>OPEN, D=>
      nx916, CLK=>clk);
   ix917 : ao32 port map ( Y=>nx916, A0=>rst, A1=>nx88, A2=>nx1325, B0=>
      signature_24_EXMPLR, B1=>nx1315);
   ix1246 : xnor2 port map ( Y=>nx1245, A0=>mult_result(24), A1=>
      signature_25_EXMPLR);
   reg_MISR_REG_25 : dff port map ( Q=>signature_25_EXMPLR, QB=>OPEN, D=>
      nx906, CLK=>clk);
   ix907 : ao32 port map ( Y=>nx906, A0=>rst, A1=>nx76, A2=>nx1325, B0=>
      signature_25_EXMPLR, B1=>nx1315);
   ix1251 : xnor2 port map ( Y=>nx1250, A0=>mult_result(25), A1=>
      signature_26_EXMPLR);
   reg_MISR_REG_26 : dff port map ( Q=>signature_26_EXMPLR, QB=>OPEN, D=>
      nx896, CLK=>clk);
   ix897 : ao32 port map ( Y=>nx896, A0=>rst, A1=>nx64, A2=>nx1325, B0=>
      signature_26_EXMPLR, B1=>nx1315);
   ix65 : xor2 port map ( Y=>nx64, A0=>mult_result(26), A1=>
      signature_27_EXMPLR);
   reg_MISR_REG_27 : dff port map ( Q=>signature_27_EXMPLR, QB=>OPEN, D=>
      nx886, CLK=>clk);
   ix887 : ao32 port map ( Y=>nx886, A0=>rst, A1=>nx54, A2=>nx1325, B0=>
      signature_27_EXMPLR, B1=>nx1315);
   ix55 : xor2 port map ( Y=>nx54, A0=>mult_result(27), A1=>
      signature_28_EXMPLR);
   reg_MISR_REG_28 : dff port map ( Q=>signature_28_EXMPLR, QB=>OPEN, D=>
      nx876, CLK=>clk);
   ix877 : ao32 port map ( Y=>nx876, A0=>rst, A1=>nx44, A2=>nx1325, B0=>
      signature_28_EXMPLR, B1=>nx1315);
   ix45 : xor2 port map ( Y=>nx44, A0=>mult_result(28), A1=>
      signature_29_EXMPLR);
   reg_MISR_REG_29 : dff port map ( Q=>signature_29_EXMPLR, QB=>OPEN, D=>
      nx866, CLK=>clk);
   ix867 : ao32 port map ( Y=>nx866, A0=>rst, A1=>nx34, A2=>nx1325, B0=>
      signature_29_EXMPLR, B1=>nx1315);
   ix1265 : xnor2 port map ( Y=>nx1264, A0=>mult_result(29), A1=>
      signature_30_EXMPLR);
   reg_MISR_REG_30 : dff port map ( Q=>signature_30_EXMPLR, QB=>OPEN, D=>
      nx856, CLK=>clk);
   ix857 : ao32 port map ( Y=>nx856, A0=>rst, A1=>nx22, A2=>nx1325, B0=>
      signature_30_EXMPLR, B1=>nx1315);
   ix23 : xor2 port map ( Y=>nx22, A0=>mult_result(30), A1=>
      signature_31_EXMPLR);
   reg_MISR_REG_31 : dff port map ( Q=>signature_31_EXMPLR, QB=>OPEN, D=>
      nx846, CLK=>clk);
   ix847 : ao32 port map ( Y=>nx846, A0=>rst, A1=>nx12, A2=>nx1325, B0=>
      signature_31_EXMPLR, B1=>nx1315);
   ix837 : mux21 port map ( Y=>nx836, A0=>signature_0_EXMPLR, A1=>zeroth_in, 
      S0=>nx1276);
   reg_zeroth_in : dff port map ( Q=>zeroth_in, QB=>nx1272, D=>nx836, CLK=>
      clk);
   ix1277 : nand02 port map ( Y=>nx1276, A0=>nx1325, A1=>rst);
   ix1169 : nor02ii port map ( Y=>nx1168, A0=>nx1329, A1=>rst);
   ix89 : xor2 port map ( Y=>nx88, A0=>nx1245, A1=>nx1272);
   ix77 : xor2 port map ( Y=>nx76, A0=>nx1250, A1=>nx1272);
   ix35 : xor2 port map ( Y=>nx34, A0=>nx1264, A1=>nx1272);
   ix13 : xor2 port map ( Y=>nx12, A0=>mult_result(31), A1=>zeroth_in);
   ix1314 : nor02ii port map ( Y=>nx1315, A0=>nx1329, A1=>rst);
   ix1316 : nor02ii port map ( Y=>nx1317, A0=>nx1329, A1=>rst);
   ix1322 : inv01 port map ( Y=>nx1323, A=>enable);
   ix1324 : inv01 port map ( Y=>nx1325, A=>nx1323);
   ix1326 : inv01 port map ( Y=>nx1327, A=>nx1323);
   ix1328 : inv01 port map ( Y=>nx1329, A=>nx1323);
end Behavioral ;

library IEEE;
library gdk;
use gdk.gdk_comps.all;
use IEEE.STD_LOGIC_1164.all;

entity MAC is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      test_mode : IN std_logic ;
      Result_OUT : OUT std_logic_vector (31 DOWNTO 0)) ;
end MAC ;

architecture structural of MAC is
   component Multiplier_32
      port (
         A : IN std_logic_vector (15 DOWNTO 0) ;
         B : IN std_logic_vector (15 DOWNTO 0) ;
         Product : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   component RCFA_32
      port (
         A : IN std_logic_vector (31 DOWNTO 0) ;
         B : IN std_logic_vector (31 DOWNTO 0) ;
         Cin : IN std_logic ;
         Sum : OUT std_logic_vector (31 DOWNTO 0) ;
         Cout : OUT std_logic) ;
   end component ;
   component RegisterN_32
      port (
         clk : IN std_logic ;
         reset : IN std_logic ;
         enable : IN std_logic ;
         input : IN std_logic_vector (31 DOWNTO 0) ;
         output : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   component LFSR
      port (
         clk : IN std_logic ;
         rst : IN std_logic ;
         enable : IN std_logic ;
         bit_pattern : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   component MISR
      port (
         clk : IN std_logic ;
         rst : IN std_logic ;
         enable : IN std_logic ;
         mult_result : IN std_logic_vector (31 DOWNTO 0) ;
         signature : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   signal MultIn1_15, MultIn1_14, MultIn1_13, MultIn1_12, MultIn1_11, 
      MultIn1_10, MultIn1_9, MultIn1_8, MultIn1_7, MultIn1_6, MultIn1_5, 
      MultIn1_4, MultIn1_3, MultIn1_2, MultIn1_1, MultIn1_0, MultIn2_15, 
      MultIn2_14, MultIn2_13, MultIn2_12, MultIn2_11, MultIn2_10, MultIn2_9, 
      MultIn2_8, MultIn2_7, MultIn2_6, MultIn2_5, MultIn2_4, MultIn2_3, 
      MultIn2_2, MultIn2_1, MultIn2_0, LFSR_OUT_31, LFSR_OUT_30, LFSR_OUT_29, 
      LFSR_OUT_28, LFSR_OUT_27, LFSR_OUT_26, LFSR_OUT_25, LFSR_OUT_24, 
      LFSR_OUT_23, LFSR_OUT_22, LFSR_OUT_21, LFSR_OUT_20, LFSR_OUT_19, 
      LFSR_OUT_18, LFSR_OUT_17, LFSR_OUT_16, LFSR_OUT_15, LFSR_OUT_14, 
      LFSR_OUT_13, LFSR_OUT_12, LFSR_OUT_11, LFSR_OUT_10, LFSR_OUT_9, 
      LFSR_OUT_8, LFSR_OUT_7, LFSR_OUT_6, LFSR_OUT_5, LFSR_OUT_4, LFSR_OUT_3, 
      LFSR_OUT_2, LFSR_OUT_1, LFSR_OUT_0, MISR_OUT_31, MISR_OUT_30, 
      MISR_OUT_29, MISR_OUT_28, MISR_OUT_27, MISR_OUT_26, MISR_OUT_25, 
      MISR_OUT_24, MISR_OUT_23, MISR_OUT_22, MISR_OUT_21, MISR_OUT_20, 
      MISR_OUT_19, MISR_OUT_18, MISR_OUT_17, MISR_OUT_16, MISR_OUT_15, 
      MISR_OUT_14, MISR_OUT_13, MISR_OUT_12, MISR_OUT_11, MISR_OUT_10, 
      MISR_OUT_9, MISR_OUT_8, MISR_OUT_7, MISR_OUT_6, MISR_OUT_5, MISR_OUT_4, 
      MISR_OUT_3, MISR_OUT_2, MISR_OUT_1, MISR_OUT_0, MULT_OUT_31, 
      MULT_OUT_30, MULT_OUT_29, MULT_OUT_28, MULT_OUT_27, MULT_OUT_26, 
      MULT_OUT_25, MULT_OUT_24, MULT_OUT_23, MULT_OUT_22, MULT_OUT_21, 
      MULT_OUT_20, MULT_OUT_19, MULT_OUT_18, MULT_OUT_17, MULT_OUT_16, 
      MULT_OUT_15, MULT_OUT_14, MULT_OUT_13, MULT_OUT_12, MULT_OUT_11, 
      MULT_OUT_10, MULT_OUT_9, MULT_OUT_8, MULT_OUT_7, MULT_OUT_6, 
      MULT_OUT_5, MULT_OUT_4, MULT_OUT_3, MULT_OUT_2, MULT_OUT_1, MULT_OUT_0, 
      ADDER_OUT_31, ADDER_OUT_30, ADDER_OUT_29, ADDER_OUT_28, ADDER_OUT_27, 
      ADDER_OUT_26, ADDER_OUT_25, ADDER_OUT_24, ADDER_OUT_23, ADDER_OUT_22, 
      ADDER_OUT_21, ADDER_OUT_20, ADDER_OUT_19, ADDER_OUT_18, ADDER_OUT_17, 
      ADDER_OUT_16, ADDER_OUT_15, ADDER_OUT_14, ADDER_OUT_13, ADDER_OUT_12, 
      ADDER_OUT_11, ADDER_OUT_10, ADDER_OUT_9, ADDER_OUT_8, ADDER_OUT_7, 
      ADDER_OUT_6, ADDER_OUT_5, ADDER_OUT_4, ADDER_OUT_3, ADDER_OUT_2, 
      ADDER_OUT_1, ADDER_OUT_0, REG_OUT_31, REG_OUT_30, REG_OUT_29, 
      REG_OUT_28, REG_OUT_27, REG_OUT_26, REG_OUT_25, REG_OUT_24, REG_OUT_23, 
      REG_OUT_22, REG_OUT_21, REG_OUT_20, REG_OUT_19, REG_OUT_18, REG_OUT_17, 
      REG_OUT_16, REG_OUT_15, REG_OUT_14, REG_OUT_13, REG_OUT_12, REG_OUT_11, 
      REG_OUT_10, REG_OUT_9, REG_OUT_8, REG_OUT_7, REG_OUT_6, REG_OUT_5, 
      REG_OUT_4, REG_OUT_3, REG_OUT_2, REG_OUT_1, REG_OUT_0, MISR_EN, GND0, 
      PWR, nx0, clk_cnt_30, nx937, clk_cnt_29, clk_cnt_28, clk_cnt_27, 
      clk_cnt_26, clk_cnt_25, clk_cnt_24, clk_cnt_23, clk_cnt_22, clk_cnt_21, 
      clk_cnt_20, clk_cnt_19, clk_cnt_18, clk_cnt_17, clk_cnt_16, clk_cnt_15, 
      clk_cnt_14, clk_cnt_13, clk_cnt_12, clk_cnt_11, clk_cnt_10, clk_cnt_9, 
      clk_cnt_8, clk_cnt_7, clk_cnt_6, clk_cnt_5, clk_cnt_4, clk_cnt_3, 
      clk_cnt_2, clk_cnt_1, clk_cnt_0, nx4, nx18, nx28, nx44, nx943, nx76, 
      nx947, nx108, nx949, nx130, nx140, nx953, nx162, nx172, nx956, nx194, 
      nx204, nx959, nx226, nx236, nx963, nx258, nx268, nx965, nx290, nx300, 
      nx969, nx322, nx332, nx972, nx354, nx364, nx975, nx386, nx396, nx979, 
      nx418, nx428, nx981, nx450, nx460, nx478, nx484, nx504, nx514, nx526, 
      nx536, nx550, nx560, nx572, nx582, nx588, nx602, nx610, nx644, nx652, 
      nx662, nx991, nx1001, nx1011, nx1021, nx1031, nx1041, nx1051, nx1061, 
      nx1071, nx1081, nx1091, nx1101, nx1111, nx1121, nx1131, nx1141, nx1151, 
      nx1161, nx1171, nx1181, nx1191, nx1201, nx1211, nx1221, nx1231, nx1241, 
      nx1251, nx1261, nx1271, nx1281, nx1291, nx1299, nx1311, nx1321, nx1327, 
      nx1331, nx1334, nx1336, nx1340, nx1344, nx1347, nx1351, nx1353, nx1357, 
      nx1361, nx1364, nx1368, nx1370, nx1374, nx1378, nx1381, nx1385, nx1387, 
      nx1391, nx1395, nx1398, nx1402, nx1404, nx1408, nx1412, nx1415, nx1419, 
      nx1421, nx1425, nx1429, nx1432, nx1436, nx1438, nx1442, nx1446, nx1449, 
      nx1453, nx1455, nx1459, nx1463, nx1466, nx1470, nx1472, nx1476, nx1480, 
      nx1483, nx1487, nx1489, nx1493, nx1497, nx1500, nx1504, nx1506, nx1510, 
      nx1514, nx1517, nx1521, nx1523, nx1527, nx1530, nx1533, nx1537, nx1539, 
      nx1543, nx1546, nx1549, nx1553, nx1555, nx1558, nx1562, nx1564, nx1567, 
      nx1572, nx1590, nx1592, nx1597, nx1603, nx1608, nx1615, nx1691, nx1693, 
      nx1695, nx1697, nx1699, nx1701, nx1705, nx1711, nx1713, nx1715, nx1717, 
      nx1719, nx1721: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   Multiplier0 : Multiplier_32 port map ( A(15)=>MultIn1_15, A(14)=>
      MultIn1_14, A(13)=>MultIn1_13, A(12)=>MultIn1_12, A(11)=>MultIn1_11, 
      A(10)=>MultIn1_10, A(9)=>MultIn1_9, A(8)=>MultIn1_8, A(7)=>MultIn1_7, 
      A(6)=>MultIn1_6, A(5)=>MultIn1_5, A(4)=>MultIn1_4, A(3)=>MultIn1_3, 
      A(2)=>MultIn1_2, A(1)=>MultIn1_1, A(0)=>MultIn1_0, B(15)=>MultIn2_15, 
      B(14)=>MultIn2_14, B(13)=>MultIn2_13, B(12)=>MultIn2_12, B(11)=>
      MultIn2_11, B(10)=>MultIn2_10, B(9)=>MultIn2_9, B(8)=>MultIn2_8, B(7)
      =>MultIn2_7, B(6)=>MultIn2_6, B(5)=>MultIn2_5, B(4)=>MultIn2_4, B(3)=>
      MultIn2_3, B(2)=>MultIn2_2, B(1)=>MultIn2_1, B(0)=>MultIn2_0, 
      Product(31)=>MULT_OUT_31, Product(30)=>MULT_OUT_30, Product(29)=>
      MULT_OUT_29, Product(28)=>MULT_OUT_28, Product(27)=>MULT_OUT_27, 
      Product(26)=>MULT_OUT_26, Product(25)=>MULT_OUT_25, Product(24)=>
      MULT_OUT_24, Product(23)=>MULT_OUT_23, Product(22)=>MULT_OUT_22, 
      Product(21)=>MULT_OUT_21, Product(20)=>MULT_OUT_20, Product(19)=>
      MULT_OUT_19, Product(18)=>MULT_OUT_18, Product(17)=>MULT_OUT_17, 
      Product(16)=>MULT_OUT_16, Product(15)=>MULT_OUT_15, Product(14)=>
      MULT_OUT_14, Product(13)=>MULT_OUT_13, Product(12)=>MULT_OUT_12, 
      Product(11)=>MULT_OUT_11, Product(10)=>MULT_OUT_10, Product(9)=>
      MULT_OUT_9, Product(8)=>MULT_OUT_8, Product(7)=>MULT_OUT_7, Product(6)
      =>MULT_OUT_6, Product(5)=>MULT_OUT_5, Product(4)=>MULT_OUT_4, 
      Product(3)=>MULT_OUT_3, Product(2)=>MULT_OUT_2, Product(1)=>MULT_OUT_1, 
      Product(0)=>MULT_OUT_0);
   RCFA0 : RCFA_32 port map ( A(31)=>MULT_OUT_31, A(30)=>MULT_OUT_30, A(29)
      =>MULT_OUT_29, A(28)=>MULT_OUT_28, A(27)=>MULT_OUT_27, A(26)=>
      MULT_OUT_26, A(25)=>MULT_OUT_25, A(24)=>MULT_OUT_24, A(23)=>
      MULT_OUT_23, A(22)=>MULT_OUT_22, A(21)=>MULT_OUT_21, A(20)=>
      MULT_OUT_20, A(19)=>MULT_OUT_19, A(18)=>MULT_OUT_18, A(17)=>
      MULT_OUT_17, A(16)=>MULT_OUT_16, A(15)=>MULT_OUT_15, A(14)=>
      MULT_OUT_14, A(13)=>MULT_OUT_13, A(12)=>MULT_OUT_12, A(11)=>
      MULT_OUT_11, A(10)=>MULT_OUT_10, A(9)=>MULT_OUT_9, A(8)=>MULT_OUT_8, 
      A(7)=>MULT_OUT_7, A(6)=>MULT_OUT_6, A(5)=>MULT_OUT_5, A(4)=>MULT_OUT_4, 
      A(3)=>MULT_OUT_3, A(2)=>MULT_OUT_2, A(1)=>MULT_OUT_1, A(0)=>MULT_OUT_0, 
      B(31)=>REG_OUT_31, B(30)=>REG_OUT_30, B(29)=>REG_OUT_29, B(28)=>
      REG_OUT_28, B(27)=>REG_OUT_27, B(26)=>REG_OUT_26, B(25)=>REG_OUT_25, 
      B(24)=>REG_OUT_24, B(23)=>REG_OUT_23, B(22)=>REG_OUT_22, B(21)=>
      REG_OUT_21, B(20)=>REG_OUT_20, B(19)=>REG_OUT_19, B(18)=>REG_OUT_18, 
      B(17)=>REG_OUT_17, B(16)=>REG_OUT_16, B(15)=>REG_OUT_15, B(14)=>
      REG_OUT_14, B(13)=>REG_OUT_13, B(12)=>REG_OUT_12, B(11)=>REG_OUT_11, 
      B(10)=>REG_OUT_10, B(9)=>REG_OUT_9, B(8)=>REG_OUT_8, B(7)=>REG_OUT_7, 
      B(6)=>REG_OUT_6, B(5)=>REG_OUT_5, B(4)=>REG_OUT_4, B(3)=>REG_OUT_3, 
      B(2)=>REG_OUT_2, B(1)=>REG_OUT_1, B(0)=>REG_OUT_0, Cin=>GND0, Sum(31)
      =>ADDER_OUT_31, Sum(30)=>ADDER_OUT_30, Sum(29)=>ADDER_OUT_29, Sum(28)
      =>ADDER_OUT_28, Sum(27)=>ADDER_OUT_27, Sum(26)=>ADDER_OUT_26, Sum(25)
      =>ADDER_OUT_25, Sum(24)=>ADDER_OUT_24, Sum(23)=>ADDER_OUT_23, Sum(22)
      =>ADDER_OUT_22, Sum(21)=>ADDER_OUT_21, Sum(20)=>ADDER_OUT_20, Sum(19)
      =>ADDER_OUT_19, Sum(18)=>ADDER_OUT_18, Sum(17)=>ADDER_OUT_17, Sum(16)
      =>ADDER_OUT_16, Sum(15)=>ADDER_OUT_15, Sum(14)=>ADDER_OUT_14, Sum(13)
      =>ADDER_OUT_13, Sum(12)=>ADDER_OUT_12, Sum(11)=>ADDER_OUT_11, Sum(10)
      =>ADDER_OUT_10, Sum(9)=>ADDER_OUT_9, Sum(8)=>ADDER_OUT_8, Sum(7)=>
      ADDER_OUT_7, Sum(6)=>ADDER_OUT_6, Sum(5)=>ADDER_OUT_5, Sum(4)=>
      ADDER_OUT_4, Sum(3)=>ADDER_OUT_3, Sum(2)=>ADDER_OUT_2, Sum(1)=>
      ADDER_OUT_1, Sum(0)=>ADDER_OUT_0, Cout=>DANGLING(0));
   RegisterN0 : RegisterN_32 port map ( clk=>clk, reset=>rst, enable=>PWR, 
      input(31)=>ADDER_OUT_31, input(30)=>ADDER_OUT_30, input(29)=>
      ADDER_OUT_29, input(28)=>ADDER_OUT_28, input(27)=>ADDER_OUT_27, 
      input(26)=>ADDER_OUT_26, input(25)=>ADDER_OUT_25, input(24)=>
      ADDER_OUT_24, input(23)=>ADDER_OUT_23, input(22)=>ADDER_OUT_22, 
      input(21)=>ADDER_OUT_21, input(20)=>ADDER_OUT_20, input(19)=>
      ADDER_OUT_19, input(18)=>ADDER_OUT_18, input(17)=>ADDER_OUT_17, 
      input(16)=>ADDER_OUT_16, input(15)=>ADDER_OUT_15, input(14)=>
      ADDER_OUT_14, input(13)=>ADDER_OUT_13, input(12)=>ADDER_OUT_12, 
      input(11)=>ADDER_OUT_11, input(10)=>ADDER_OUT_10, input(9)=>
      ADDER_OUT_9, input(8)=>ADDER_OUT_8, input(7)=>ADDER_OUT_7, input(6)=>
      ADDER_OUT_6, input(5)=>ADDER_OUT_5, input(4)=>ADDER_OUT_4, input(3)=>
      ADDER_OUT_3, input(2)=>ADDER_OUT_2, input(1)=>ADDER_OUT_1, input(0)=>
      ADDER_OUT_0, output(31)=>REG_OUT_31, output(30)=>REG_OUT_30, 
      output(29)=>REG_OUT_29, output(28)=>REG_OUT_28, output(27)=>REG_OUT_27, 
      output(26)=>REG_OUT_26, output(25)=>REG_OUT_25, output(24)=>REG_OUT_24, 
      output(23)=>REG_OUT_23, output(22)=>REG_OUT_22, output(21)=>REG_OUT_21, 
      output(20)=>REG_OUT_20, output(19)=>REG_OUT_19, output(18)=>REG_OUT_18, 
      output(17)=>REG_OUT_17, output(16)=>REG_OUT_16, output(15)=>REG_OUT_15, 
      output(14)=>REG_OUT_14, output(13)=>REG_OUT_13, output(12)=>REG_OUT_12, 
      output(11)=>REG_OUT_11, output(10)=>REG_OUT_10, output(9)=>REG_OUT_9, 
      output(8)=>REG_OUT_8, output(7)=>REG_OUT_7, output(6)=>REG_OUT_6, 
      output(5)=>REG_OUT_5, output(4)=>REG_OUT_4, output(3)=>REG_OUT_3, 
      output(2)=>REG_OUT_2, output(1)=>REG_OUT_1, output(0)=>REG_OUT_0);
   LFSR0 : LFSR port map ( clk=>clk, rst=>rst, enable=>test_mode, 
      bit_pattern(31)=>LFSR_OUT_31, bit_pattern(30)=>LFSR_OUT_30, 
      bit_pattern(29)=>LFSR_OUT_29, bit_pattern(28)=>LFSR_OUT_28, 
      bit_pattern(27)=>LFSR_OUT_27, bit_pattern(26)=>LFSR_OUT_26, 
      bit_pattern(25)=>LFSR_OUT_25, bit_pattern(24)=>LFSR_OUT_24, 
      bit_pattern(23)=>LFSR_OUT_23, bit_pattern(22)=>LFSR_OUT_22, 
      bit_pattern(21)=>LFSR_OUT_21, bit_pattern(20)=>LFSR_OUT_20, 
      bit_pattern(19)=>LFSR_OUT_19, bit_pattern(18)=>LFSR_OUT_18, 
      bit_pattern(17)=>LFSR_OUT_17, bit_pattern(16)=>LFSR_OUT_16, 
      bit_pattern(15)=>LFSR_OUT_15, bit_pattern(14)=>LFSR_OUT_14, 
      bit_pattern(13)=>LFSR_OUT_13, bit_pattern(12)=>LFSR_OUT_12, 
      bit_pattern(11)=>LFSR_OUT_11, bit_pattern(10)=>LFSR_OUT_10, 
      bit_pattern(9)=>LFSR_OUT_9, bit_pattern(8)=>LFSR_OUT_8, bit_pattern(7)
      =>LFSR_OUT_7, bit_pattern(6)=>LFSR_OUT_6, bit_pattern(5)=>LFSR_OUT_5, 
      bit_pattern(4)=>LFSR_OUT_4, bit_pattern(3)=>LFSR_OUT_3, bit_pattern(2)
      =>LFSR_OUT_2, bit_pattern(1)=>LFSR_OUT_1, bit_pattern(0)=>LFSR_OUT_0);
   MISR0 : MISR port map ( clk=>clk, rst=>rst, enable=>MISR_EN, 
      mult_result(31)=>REG_OUT_31, mult_result(30)=>REG_OUT_30, 
      mult_result(29)=>REG_OUT_29, mult_result(28)=>REG_OUT_28, 
      mult_result(27)=>REG_OUT_27, mult_result(26)=>REG_OUT_26, 
      mult_result(25)=>REG_OUT_25, mult_result(24)=>REG_OUT_24, 
      mult_result(23)=>REG_OUT_23, mult_result(22)=>REG_OUT_22, 
      mult_result(21)=>REG_OUT_21, mult_result(20)=>REG_OUT_20, 
      mult_result(19)=>REG_OUT_19, mult_result(18)=>REG_OUT_18, 
      mult_result(17)=>REG_OUT_17, mult_result(16)=>REG_OUT_16, 
      mult_result(15)=>REG_OUT_15, mult_result(14)=>REG_OUT_14, 
      mult_result(13)=>REG_OUT_13, mult_result(12)=>REG_OUT_12, 
      mult_result(11)=>REG_OUT_11, mult_result(10)=>REG_OUT_10, 
      mult_result(9)=>REG_OUT_9, mult_result(8)=>REG_OUT_8, mult_result(7)=>
      REG_OUT_7, mult_result(6)=>REG_OUT_6, mult_result(5)=>REG_OUT_5, 
      mult_result(4)=>REG_OUT_4, mult_result(3)=>REG_OUT_3, mult_result(2)=>
      REG_OUT_2, mult_result(1)=>REG_OUT_1, mult_result(0)=>REG_OUT_0, 
      signature(31)=>MISR_OUT_31, signature(30)=>MISR_OUT_30, signature(29)
      =>MISR_OUT_29, signature(28)=>MISR_OUT_28, signature(27)=>MISR_OUT_27, 
      signature(26)=>MISR_OUT_26, signature(25)=>MISR_OUT_25, signature(24)
      =>MISR_OUT_24, signature(23)=>MISR_OUT_23, signature(22)=>MISR_OUT_22, 
      signature(21)=>MISR_OUT_21, signature(20)=>MISR_OUT_20, signature(19)
      =>MISR_OUT_19, signature(18)=>MISR_OUT_18, signature(17)=>MISR_OUT_17, 
      signature(16)=>MISR_OUT_16, signature(15)=>MISR_OUT_15, signature(14)
      =>MISR_OUT_14, signature(13)=>MISR_OUT_13, signature(12)=>MISR_OUT_12, 
      signature(11)=>MISR_OUT_11, signature(10)=>MISR_OUT_10, signature(9)=>
      MISR_OUT_9, signature(8)=>MISR_OUT_8, signature(7)=>MISR_OUT_7, 
      signature(6)=>MISR_OUT_6, signature(5)=>MISR_OUT_5, signature(4)=>
      MISR_OUT_4, signature(3)=>MISR_OUT_3, signature(2)=>MISR_OUT_2, 
      signature(1)=>MISR_OUT_1, signature(0)=>MISR_OUT_0);
   ix799 : fake_vcc port map ( Y=>PWR);
   ix797 : fake_gnd port map ( Y=>GND0);
   reg_MISR_EN : dff port map ( Q=>MISR_EN, QB=>OPEN, D=>nx1311, CLK=>clk);
   ix663 : mux21 port map ( Y=>nx662, A0=>MISR_EN, A1=>nx610, S0=>nx1615);
   ix611 : oai21 port map ( Y=>nx610, A0=>nx1321, A1=>nx1597, B0=>nx1608);
   ix1322 : nand04 port map ( Y=>nx1321, A0=>nx504, A1=>nx514, A2=>nx526, A3
      =>nx536);
   ix485 : aoi21 port map ( Y=>nx484, A0=>nx1327, A1=>nx1590, B0=>nx1592);
   ix1328 : nand02 port map ( Y=>nx1327, A0=>clk_cnt_29, A1=>nx981);
   ix1282 : oai21 port map ( Y=>nx1281, A0=>nx1331, A1=>nx1693, B0=>nx1336);
   reg_clk_cnt_29 : dff port map ( Q=>clk_cnt_29, QB=>nx1331, D=>nx1281, CLK
      =>clk);
   ix1335 : nand02 port map ( Y=>nx1334, A0=>rst, A1=>test_mode);
   ix1337 : nand04 port map ( Y=>nx1336, A0=>nx460, A1=>nx0, A2=>nx1327, A3
      =>nx1697);
   ix461 : or02 port map ( Y=>nx460, A0=>nx981, A1=>clk_cnt_29);
   ix451 : nor03 port map ( Y=>nx450, A0=>nx1344, A1=>nx1699, A2=>nx981);
   reg_clk_cnt_28 : dff port map ( Q=>clk_cnt_28, QB=>nx1340, D=>nx1271, CLK
      =>clk);
   ix1348 : nand02 port map ( Y=>nx1347, A0=>clk_cnt_27, A1=>nx979);
   ix1262 : oai21 port map ( Y=>nx1261, A0=>nx1351, A1=>nx1693, B0=>nx1353);
   reg_clk_cnt_27 : dff port map ( Q=>clk_cnt_27, QB=>nx1351, D=>nx1261, CLK
      =>clk);
   ix1354 : nand04 port map ( Y=>nx1353, A0=>nx428, A1=>nx0, A2=>nx1347, A3
      =>nx1697);
   ix429 : or02 port map ( Y=>nx428, A0=>nx979, A1=>clk_cnt_27);
   ix419 : nor03 port map ( Y=>nx418, A0=>nx1361, A1=>nx1699, A2=>nx979);
   reg_clk_cnt_26 : dff port map ( Q=>clk_cnt_26, QB=>nx1357, D=>nx1251, CLK
      =>clk);
   ix1365 : nand02 port map ( Y=>nx1364, A0=>clk_cnt_25, A1=>nx975);
   ix1242 : oai21 port map ( Y=>nx1241, A0=>nx1368, A1=>nx1693, B0=>nx1370);
   reg_clk_cnt_25 : dff port map ( Q=>clk_cnt_25, QB=>nx1368, D=>nx1241, CLK
      =>clk);
   ix1371 : nand04 port map ( Y=>nx1370, A0=>nx396, A1=>nx0, A2=>nx1364, A3
      =>nx1697);
   ix397 : or02 port map ( Y=>nx396, A0=>nx975, A1=>clk_cnt_25);
   ix387 : nor03 port map ( Y=>nx386, A0=>nx1378, A1=>nx1699, A2=>nx975);
   reg_clk_cnt_24 : dff port map ( Q=>clk_cnt_24, QB=>nx1374, D=>nx1231, CLK
      =>clk);
   ix1382 : nand02 port map ( Y=>nx1381, A0=>clk_cnt_23, A1=>nx972);
   ix1222 : oai21 port map ( Y=>nx1221, A0=>nx1385, A1=>nx1693, B0=>nx1387);
   reg_clk_cnt_23 : dff port map ( Q=>clk_cnt_23, QB=>nx1385, D=>nx1221, CLK
      =>clk);
   ix1388 : nand04 port map ( Y=>nx1387, A0=>nx364, A1=>nx0, A2=>nx1381, A3
      =>nx1697);
   ix365 : or02 port map ( Y=>nx364, A0=>nx972, A1=>clk_cnt_23);
   ix355 : nor03 port map ( Y=>nx354, A0=>nx1395, A1=>nx1699, A2=>nx972);
   reg_clk_cnt_22 : dff port map ( Q=>clk_cnt_22, QB=>nx1391, D=>nx1211, CLK
      =>clk);
   ix1399 : nand02 port map ( Y=>nx1398, A0=>clk_cnt_21, A1=>nx969);
   ix1202 : oai21 port map ( Y=>nx1201, A0=>nx1402, A1=>nx1693, B0=>nx1404);
   reg_clk_cnt_21 : dff port map ( Q=>clk_cnt_21, QB=>nx1402, D=>nx1201, CLK
      =>clk);
   ix1405 : nand04 port map ( Y=>nx1404, A0=>nx332, A1=>nx1691, A2=>nx1398, 
      A3=>nx1695);
   ix333 : or02 port map ( Y=>nx332, A0=>nx969, A1=>clk_cnt_21);
   ix323 : nor03 port map ( Y=>nx322, A0=>nx1412, A1=>nx1699, A2=>nx969);
   reg_clk_cnt_20 : dff port map ( Q=>clk_cnt_20, QB=>nx1408, D=>nx1191, CLK
      =>clk);
   ix1416 : nand02 port map ( Y=>nx1415, A0=>clk_cnt_19, A1=>nx965);
   ix1182 : oai21 port map ( Y=>nx1181, A0=>nx1419, A1=>nx1693, B0=>nx1421);
   reg_clk_cnt_19 : dff port map ( Q=>clk_cnt_19, QB=>nx1419, D=>nx1181, CLK
      =>clk);
   ix1422 : nand04 port map ( Y=>nx1421, A0=>nx300, A1=>nx1691, A2=>nx1415, 
      A3=>nx1695);
   ix301 : or02 port map ( Y=>nx300, A0=>nx965, A1=>clk_cnt_19);
   ix291 : nor03 port map ( Y=>nx290, A0=>nx1429, A1=>nx1699, A2=>nx965);
   reg_clk_cnt_18 : dff port map ( Q=>clk_cnt_18, QB=>nx1425, D=>nx1171, CLK
      =>clk);
   ix1433 : nand02 port map ( Y=>nx1432, A0=>clk_cnt_17, A1=>nx963);
   ix1162 : oai21 port map ( Y=>nx1161, A0=>nx1436, A1=>nx1693, B0=>nx1438);
   reg_clk_cnt_17 : dff port map ( Q=>clk_cnt_17, QB=>nx1436, D=>nx1161, CLK
      =>clk);
   ix1439 : nand04 port map ( Y=>nx1438, A0=>nx268, A1=>nx1691, A2=>nx1432, 
      A3=>nx1695);
   ix269 : or02 port map ( Y=>nx268, A0=>nx963, A1=>clk_cnt_17);
   ix259 : nor03 port map ( Y=>nx258, A0=>nx1446, A1=>nx1699, A2=>nx963);
   reg_clk_cnt_16 : dff port map ( Q=>clk_cnt_16, QB=>nx1442, D=>nx1151, CLK
      =>clk);
   ix1450 : nand02 port map ( Y=>nx1449, A0=>clk_cnt_15, A1=>nx959);
   ix1142 : oai21 port map ( Y=>nx1141, A0=>nx1453, A1=>nx1693, B0=>nx1455);
   reg_clk_cnt_15 : dff port map ( Q=>clk_cnt_15, QB=>nx1453, D=>nx1141, CLK
      =>clk);
   ix1456 : nand04 port map ( Y=>nx1455, A0=>nx236, A1=>nx1691, A2=>nx1449, 
      A3=>nx1695);
   ix237 : or02 port map ( Y=>nx236, A0=>nx959, A1=>clk_cnt_15);
   ix227 : nor03 port map ( Y=>nx226, A0=>nx1463, A1=>nx1699, A2=>nx959);
   reg_clk_cnt_14 : dff port map ( Q=>clk_cnt_14, QB=>nx1459, D=>nx1131, CLK
      =>clk);
   ix1467 : nand02 port map ( Y=>nx1466, A0=>clk_cnt_13, A1=>nx956);
   ix1122 : oai21 port map ( Y=>nx1121, A0=>nx1470, A1=>nx1693, B0=>nx1472);
   reg_clk_cnt_13 : dff port map ( Q=>clk_cnt_13, QB=>nx1470, D=>nx1121, CLK
      =>clk);
   ix1473 : nand04 port map ( Y=>nx1472, A0=>nx204, A1=>nx1691, A2=>nx1466, 
      A3=>nx1695);
   ix205 : or02 port map ( Y=>nx204, A0=>nx956, A1=>clk_cnt_13);
   ix195 : nor03 port map ( Y=>nx194, A0=>nx1480, A1=>nx1699, A2=>nx956);
   reg_clk_cnt_12 : dff port map ( Q=>clk_cnt_12, QB=>nx1476, D=>nx1111, CLK
      =>clk);
   ix1484 : nand02 port map ( Y=>nx1483, A0=>clk_cnt_11, A1=>nx953);
   ix1102 : oai21 port map ( Y=>nx1101, A0=>nx1487, A1=>nx1693, B0=>nx1489);
   reg_clk_cnt_11 : dff port map ( Q=>clk_cnt_11, QB=>nx1487, D=>nx1101, CLK
      =>clk);
   ix1490 : nand04 port map ( Y=>nx1489, A0=>nx172, A1=>nx1691, A2=>nx1483, 
      A3=>nx1695);
   ix173 : or02 port map ( Y=>nx172, A0=>nx953, A1=>clk_cnt_11);
   ix163 : nor03 port map ( Y=>nx162, A0=>nx1497, A1=>nx1699, A2=>nx953);
   reg_clk_cnt_10 : dff port map ( Q=>clk_cnt_10, QB=>nx1493, D=>nx1091, CLK
      =>clk);
   ix1501 : nand02 port map ( Y=>nx1500, A0=>clk_cnt_9, A1=>nx949);
   ix1082 : oai21 port map ( Y=>nx1081, A0=>nx1504, A1=>nx1693, B0=>nx1506);
   reg_clk_cnt_9 : dff port map ( Q=>clk_cnt_9, QB=>nx1504, D=>nx1081, CLK=>
      clk);
   ix1507 : nand04 port map ( Y=>nx1506, A0=>nx140, A1=>nx1691, A2=>nx1500, 
      A3=>nx1695);
   ix141 : or02 port map ( Y=>nx140, A0=>nx949, A1=>clk_cnt_9);
   ix131 : nor03 port map ( Y=>nx130, A0=>nx1514, A1=>nx1699, A2=>nx949);
   reg_clk_cnt_8 : dff port map ( Q=>clk_cnt_8, QB=>nx1510, D=>nx1071, CLK=>
      clk);
   ix1518 : nand02 port map ( Y=>nx1517, A0=>clk_cnt_7, A1=>nx947);
   ix1062 : oai21 port map ( Y=>nx1061, A0=>nx1521, A1=>nx1693, B0=>nx1523);
   reg_clk_cnt_7 : dff port map ( Q=>clk_cnt_7, QB=>nx1521, D=>nx1061, CLK=>
      clk);
   ix1524 : nand04 port map ( Y=>nx1523, A0=>nx108, A1=>nx1691, A2=>nx1517, 
      A3=>nx1695);
   ix109 : or02 port map ( Y=>nx108, A0=>nx947, A1=>clk_cnt_7);
   ix1052 : oai21 port map ( Y=>nx1051, A0=>nx1527, A1=>nx1693, B0=>nx1530);
   ix1534 : nand02 port map ( Y=>nx1533, A0=>clk_cnt_5, A1=>nx943);
   ix1042 : oai21 port map ( Y=>nx1041, A0=>nx1537, A1=>nx1693, B0=>nx1539);
   reg_clk_cnt_5 : dff port map ( Q=>clk_cnt_5, QB=>nx1537, D=>nx1041, CLK=>
      clk);
   ix1540 : nand04 port map ( Y=>nx1539, A0=>nx76, A1=>nx1691, A2=>nx1533, 
      A3=>nx1695);
   ix77 : or02 port map ( Y=>nx76, A0=>nx943, A1=>clk_cnt_5);
   ix1032 : oai21 port map ( Y=>nx1031, A0=>nx1543, A1=>nx1693, B0=>nx1546);
   ix1550 : nand04 port map ( Y=>nx1549, A0=>clk_cnt_3, A1=>clk_cnt_2, A2=>
      clk_cnt_1, A3=>clk_cnt_0);
   ix1022 : oai21 port map ( Y=>nx1021, A0=>nx1553, A1=>nx1695, B0=>nx1555);
   reg_clk_cnt_3 : dff port map ( Q=>clk_cnt_3, QB=>nx1553, D=>nx1021, CLK=>
      clk);
   ix1556 : nand04 port map ( Y=>nx1555, A0=>nx44, A1=>nx1691, A2=>nx1549, 
      A3=>nx1695);
   ix45 : nand02 port map ( Y=>nx44, A0=>nx1558, A1=>nx1553);
   ix1559 : nand03 port map ( Y=>nx1558, A0=>clk_cnt_2, A1=>clk_cnt_1, A2=>
      clk_cnt_0);
   ix1012 : oai21 port map ( Y=>nx1011, A0=>nx1562, A1=>nx1695, B0=>nx1564);
   reg_clk_cnt_2 : dff port map ( Q=>clk_cnt_2, QB=>nx1562, D=>nx1011, CLK=>
      clk);
   ix1565 : nand04 port map ( Y=>nx1564, A0=>nx28, A1=>nx1691, A2=>nx1558, 
      A3=>nx1695);
   ix29 : nand02 port map ( Y=>nx28, A0=>nx1567, A1=>nx1562);
   ix1568 : nand02 port map ( Y=>nx1567, A0=>clk_cnt_1, A1=>clk_cnt_0);
   reg_clk_cnt_1 : dff port map ( Q=>clk_cnt_1, QB=>OPEN, D=>nx1001, CLK=>
      clk);
   ix1573 : oai21 port map ( Y=>nx1572, A0=>clk_cnt_0, A1=>clk_cnt_1, B0=>
      nx1567);
   reg_clk_cnt_0 : dff port map ( Q=>clk_cnt_0, QB=>OPEN, D=>nx991, CLK=>clk
   );
   reg_clk_cnt_4 : dff port map ( Q=>clk_cnt_4, QB=>nx1543, D=>nx1031, CLK=>
      clk);
   reg_clk_cnt_6 : dff port map ( Q=>clk_cnt_6, QB=>nx1527, D=>nx1051, CLK=>
      clk);
   reg_clk_cnt_30 : dff port map ( Q=>clk_cnt_30, QB=>nx1590, D=>nx1291, CLK
      =>clk);
   ix1593 : oai21 port map ( Y=>nx1592, A0=>nx1590, A1=>nx1327, B0=>nx1691);
   ix1598 : nand04 port map ( Y=>nx1597, A0=>nx550, A1=>nx560, A2=>nx572, A3
      =>nx602);
   ix603 : nor03 port map ( Y=>nx602, A0=>nx1603, A1=>clk_cnt_8, A2=>
      clk_cnt_7);
   ix1604 : aoi21 port map ( Y=>nx1603, A0=>nx582, A1=>nx588, B0=>nx1527);
   clk_cnt_31 : dff port map ( Q=>OPEN, QB=>nx1608, D=>nx1299, CLK=>clk);
   ix645 : oai21 port map ( Y=>nx644, A0=>clk_cnt_1, A1=>clk_cnt_0, B0=>
      clk_cnt_2);
   ix805 : mux21 port map ( Y=>MultIn2_0, A0=>B(0), A1=>LFSR_OUT_0, S0=>
      test_mode);
   ix813 : mux21 port map ( Y=>MultIn2_1, A0=>B(1), A1=>LFSR_OUT_1, S0=>
      test_mode);
   ix821 : mux21 port map ( Y=>MultIn2_2, A0=>B(2), A1=>LFSR_OUT_2, S0=>
      test_mode);
   ix829 : mux21 port map ( Y=>MultIn2_3, A0=>B(3), A1=>LFSR_OUT_3, S0=>
      test_mode);
   ix837 : mux21 port map ( Y=>MultIn2_4, A0=>B(4), A1=>LFSR_OUT_4, S0=>
      test_mode);
   ix845 : mux21 port map ( Y=>MultIn2_5, A0=>B(5), A1=>LFSR_OUT_5, S0=>
      test_mode);
   ix853 : mux21 port map ( Y=>MultIn2_6, A0=>B(6), A1=>LFSR_OUT_6, S0=>
      test_mode);
   ix861 : mux21 port map ( Y=>MultIn2_7, A0=>B(7), A1=>LFSR_OUT_7, S0=>
      test_mode);
   ix869 : mux21 port map ( Y=>MultIn2_8, A0=>B(8), A1=>LFSR_OUT_8, S0=>
      test_mode);
   ix877 : mux21 port map ( Y=>MultIn2_9, A0=>B(9), A1=>LFSR_OUT_9, S0=>
      test_mode);
   ix885 : mux21 port map ( Y=>MultIn2_10, A0=>B(10), A1=>LFSR_OUT_10, S0=>
      test_mode);
   ix893 : mux21 port map ( Y=>MultIn2_11, A0=>B(11), A1=>LFSR_OUT_11, S0=>
      test_mode);
   ix901 : mux21 port map ( Y=>MultIn2_12, A0=>B(12), A1=>LFSR_OUT_12, S0=>
      test_mode);
   ix909 : mux21 port map ( Y=>MultIn2_13, A0=>B(13), A1=>LFSR_OUT_13, S0=>
      test_mode);
   ix917 : mux21 port map ( Y=>MultIn2_14, A0=>B(14), A1=>LFSR_OUT_14, S0=>
      test_mode);
   ix925 : mux21 port map ( Y=>MultIn2_15, A0=>B(15), A1=>LFSR_OUT_15, S0=>
      test_mode);
   ix677 : mux21 port map ( Y=>MultIn1_0, A0=>A(0), A1=>LFSR_OUT_16, S0=>
      test_mode);
   ix685 : mux21 port map ( Y=>MultIn1_1, A0=>A(1), A1=>LFSR_OUT_17, S0=>
      test_mode);
   ix693 : mux21 port map ( Y=>MultIn1_2, A0=>A(2), A1=>LFSR_OUT_18, S0=>
      test_mode);
   ix701 : mux21 port map ( Y=>MultIn1_3, A0=>A(3), A1=>LFSR_OUT_19, S0=>
      test_mode);
   ix709 : mux21 port map ( Y=>MultIn1_4, A0=>A(4), A1=>LFSR_OUT_20, S0=>
      test_mode);
   ix717 : mux21 port map ( Y=>MultIn1_5, A0=>A(5), A1=>LFSR_OUT_21, S0=>
      test_mode);
   ix725 : mux21 port map ( Y=>MultIn1_6, A0=>A(6), A1=>LFSR_OUT_22, S0=>
      test_mode);
   ix733 : mux21 port map ( Y=>MultIn1_7, A0=>A(7), A1=>LFSR_OUT_23, S0=>
      test_mode);
   ix741 : mux21 port map ( Y=>MultIn1_8, A0=>A(8), A1=>LFSR_OUT_24, S0=>
      test_mode);
   ix749 : mux21 port map ( Y=>MultIn1_9, A0=>A(9), A1=>LFSR_OUT_25, S0=>
      test_mode);
   ix757 : mux21 port map ( Y=>MultIn1_10, A0=>A(10), A1=>LFSR_OUT_26, S0=>
      test_mode);
   ix765 : mux21 port map ( Y=>MultIn1_11, A0=>A(11), A1=>LFSR_OUT_27, S0=>
      test_mode);
   ix773 : mux21 port map ( Y=>MultIn1_12, A0=>A(12), A1=>LFSR_OUT_28, S0=>
      test_mode);
   ix781 : mux21 port map ( Y=>MultIn1_13, A0=>A(13), A1=>LFSR_OUT_29, S0=>
      test_mode);
   ix789 : mux21 port map ( Y=>MultIn1_14, A0=>A(14), A1=>LFSR_OUT_30, S0=>
      test_mode);
   ix801 : mux21 port map ( Y=>MultIn1_15, A0=>A(15), A1=>LFSR_OUT_31, S0=>
      test_mode);
   ix933 : mux21 port map ( Y=>Result_OUT(0), A0=>REG_OUT_0, A1=>MISR_OUT_0, 
      S0=>test_mode);
   ix941 : mux21 port map ( Y=>Result_OUT(1), A0=>REG_OUT_1, A1=>MISR_OUT_1, 
      S0=>test_mode);
   ix949 : mux21 port map ( Y=>Result_OUT(2), A0=>REG_OUT_2, A1=>MISR_OUT_2, 
      S0=>test_mode);
   ix957 : mux21 port map ( Y=>Result_OUT(3), A0=>REG_OUT_3, A1=>MISR_OUT_3, 
      S0=>test_mode);
   ix965 : mux21 port map ( Y=>Result_OUT(4), A0=>REG_OUT_4, A1=>MISR_OUT_4, 
      S0=>test_mode);
   ix973 : mux21 port map ( Y=>Result_OUT(5), A0=>REG_OUT_5, A1=>MISR_OUT_5, 
      S0=>test_mode);
   ix981 : mux21 port map ( Y=>Result_OUT(6), A0=>REG_OUT_6, A1=>MISR_OUT_6, 
      S0=>test_mode);
   ix989 : mux21 port map ( Y=>Result_OUT(7), A0=>REG_OUT_7, A1=>MISR_OUT_7, 
      S0=>test_mode);
   ix997 : mux21 port map ( Y=>Result_OUT(8), A0=>REG_OUT_8, A1=>MISR_OUT_8, 
      S0=>test_mode);
   ix1005 : mux21 port map ( Y=>Result_OUT(9), A0=>REG_OUT_9, A1=>MISR_OUT_9, 
      S0=>test_mode);
   ix1013 : mux21 port map ( Y=>Result_OUT(10), A0=>REG_OUT_10, A1=>
      MISR_OUT_10, S0=>test_mode);
   ix1021 : mux21 port map ( Y=>Result_OUT(11), A0=>REG_OUT_11, A1=>
      MISR_OUT_11, S0=>test_mode);
   ix1029 : mux21 port map ( Y=>Result_OUT(12), A0=>REG_OUT_12, A1=>
      MISR_OUT_12, S0=>test_mode);
   ix1037 : mux21 port map ( Y=>Result_OUT(13), A0=>REG_OUT_13, A1=>
      MISR_OUT_13, S0=>test_mode);
   ix1045 : mux21 port map ( Y=>Result_OUT(14), A0=>REG_OUT_14, A1=>
      MISR_OUT_14, S0=>test_mode);
   ix1053 : mux21 port map ( Y=>Result_OUT(15), A0=>REG_OUT_15, A1=>
      MISR_OUT_15, S0=>test_mode);
   ix1061 : mux21 port map ( Y=>Result_OUT(16), A0=>REG_OUT_16, A1=>
      MISR_OUT_16, S0=>test_mode);
   ix1069 : mux21 port map ( Y=>Result_OUT(17), A0=>REG_OUT_17, A1=>
      MISR_OUT_17, S0=>test_mode);
   ix1077 : mux21 port map ( Y=>Result_OUT(18), A0=>REG_OUT_18, A1=>
      MISR_OUT_18, S0=>test_mode);
   ix1085 : mux21 port map ( Y=>Result_OUT(19), A0=>REG_OUT_19, A1=>
      MISR_OUT_19, S0=>test_mode);
   ix1093 : mux21 port map ( Y=>Result_OUT(20), A0=>REG_OUT_20, A1=>
      MISR_OUT_20, S0=>test_mode);
   ix1101 : mux21 port map ( Y=>Result_OUT(21), A0=>REG_OUT_21, A1=>
      MISR_OUT_21, S0=>test_mode);
   ix1109 : mux21 port map ( Y=>Result_OUT(22), A0=>REG_OUT_22, A1=>
      MISR_OUT_22, S0=>test_mode);
   ix1117 : mux21 port map ( Y=>Result_OUT(23), A0=>REG_OUT_23, A1=>
      MISR_OUT_23, S0=>test_mode);
   ix1125 : mux21 port map ( Y=>Result_OUT(24), A0=>REG_OUT_24, A1=>
      MISR_OUT_24, S0=>test_mode);
   ix1133 : mux21 port map ( Y=>Result_OUT(25), A0=>REG_OUT_25, A1=>
      MISR_OUT_25, S0=>test_mode);
   ix1141 : mux21 port map ( Y=>Result_OUT(26), A0=>REG_OUT_26, A1=>
      MISR_OUT_26, S0=>test_mode);
   ix1149 : mux21 port map ( Y=>Result_OUT(27), A0=>REG_OUT_27, A1=>
      MISR_OUT_27, S0=>test_mode);
   ix1157 : mux21 port map ( Y=>Result_OUT(28), A0=>REG_OUT_28, A1=>
      MISR_OUT_28, S0=>test_mode);
   ix1165 : mux21 port map ( Y=>Result_OUT(29), A0=>REG_OUT_29, A1=>
      MISR_OUT_29, S0=>test_mode);
   ix1173 : mux21 port map ( Y=>Result_OUT(30), A0=>REG_OUT_30, A1=>
      MISR_OUT_30, S0=>test_mode);
   ix1181 : mux21 port map ( Y=>Result_OUT(31), A0=>REG_OUT_31, A1=>
      MISR_OUT_31, S0=>test_mode);
   ix1 : inv01 port map ( Y=>nx0, A=>nx1334);
   ix1690 : inv01 port map ( Y=>nx1691, A=>nx1701);
   ix1692 : inv02 port map ( Y=>nx1693, A=>nx1705);
   ix1694 : inv02 port map ( Y=>nx1695, A=>nx1705);
   ix1696 : inv02 port map ( Y=>nx1697, A=>nx1705);
   ix1698 : inv01 port map ( Y=>nx1699, A=>nx0);
   ix1700 : inv01 port map ( Y=>nx1701, A=>nx0);
   ix1704 : inv02 port map ( Y=>nx1705, A=>nx937);
   ix1312 : mux21 port map ( Y=>nx1311, A0=>MISR_EN, A1=>nx662, S0=>nx0);
   ix505 : and04 port map ( Y=>nx504, A0=>nx1590, A1=>nx1331, A2=>nx1340, A3
      =>nx1351);
   ix1292 : mux21 port map ( Y=>nx1291, A0=>clk_cnt_30, A1=>nx484, S0=>
      nx1719);
   ix459 : nor02ii port map ( Y=>nx981, A0=>nx1347, A1=>clk_cnt_28);
   ix1272 : mux21 port map ( Y=>nx1271, A0=>clk_cnt_28, A1=>nx450, S0=>
      nx1719);
   ix1345 : and02 port map ( Y=>nx1344, A0=>nx1340, A1=>nx1347);
   ix427 : nor02ii port map ( Y=>nx979, A0=>nx1364, A1=>clk_cnt_26);
   ix1252 : mux21 port map ( Y=>nx1251, A0=>clk_cnt_26, A1=>nx418, S0=>
      nx1719);
   ix1362 : and02 port map ( Y=>nx1361, A0=>nx1357, A1=>nx1364);
   ix395 : nor02ii port map ( Y=>nx975, A0=>nx1381, A1=>clk_cnt_24);
   ix1232 : mux21 port map ( Y=>nx1231, A0=>clk_cnt_24, A1=>nx386, S0=>
      nx1719);
   ix1379 : and02 port map ( Y=>nx1378, A0=>nx1374, A1=>nx1381);
   ix363 : nor02ii port map ( Y=>nx972, A0=>nx1398, A1=>clk_cnt_22);
   ix1212 : mux21 port map ( Y=>nx1211, A0=>clk_cnt_22, A1=>nx354, S0=>
      nx1719);
   ix1396 : and02 port map ( Y=>nx1395, A0=>nx1391, A1=>nx1398);
   ix331 : nor02ii port map ( Y=>nx969, A0=>nx1415, A1=>clk_cnt_20);
   ix1192 : mux21 port map ( Y=>nx1191, A0=>clk_cnt_20, A1=>nx322, S0=>
      nx1719);
   ix1413 : and02 port map ( Y=>nx1412, A0=>nx1408, A1=>nx1415);
   ix299 : nor02ii port map ( Y=>nx965, A0=>nx1432, A1=>clk_cnt_18);
   ix1172 : mux21 port map ( Y=>nx1171, A0=>clk_cnt_18, A1=>nx290, S0=>
      nx1719);
   ix1430 : and02 port map ( Y=>nx1429, A0=>nx1425, A1=>nx1432);
   ix267 : nor02ii port map ( Y=>nx963, A0=>nx1449, A1=>clk_cnt_16);
   ix1152 : mux21 port map ( Y=>nx1151, A0=>clk_cnt_16, A1=>nx258, S0=>
      nx1719);
   ix1447 : and02 port map ( Y=>nx1446, A0=>nx1442, A1=>nx1449);
   ix235 : nor02ii port map ( Y=>nx959, A0=>nx1466, A1=>clk_cnt_14);
   ix1132 : mux21 port map ( Y=>nx1131, A0=>clk_cnt_14, A1=>nx226, S0=>
      nx1719);
   ix1464 : and02 port map ( Y=>nx1463, A0=>nx1459, A1=>nx1466);
   ix203 : nor02ii port map ( Y=>nx956, A0=>nx1483, A1=>clk_cnt_12);
   ix1112 : mux21 port map ( Y=>nx1111, A0=>clk_cnt_12, A1=>nx194, S0=>
      nx1719);
   ix1481 : and02 port map ( Y=>nx1480, A0=>nx1476, A1=>nx1483);
   ix171 : nor02ii port map ( Y=>nx953, A0=>nx1500, A1=>clk_cnt_10);
   ix1092 : mux21 port map ( Y=>nx1091, A0=>clk_cnt_10, A1=>nx162, S0=>
      nx1721);
   ix1498 : and02 port map ( Y=>nx1497, A0=>nx1493, A1=>nx1500);
   ix139 : nor02ii port map ( Y=>nx949, A0=>nx1517, A1=>clk_cnt_8);
   ix1072 : mux21 port map ( Y=>nx1071, A0=>clk_cnt_8, A1=>nx130, S0=>nx1721
   );
   ix1515 : and02 port map ( Y=>nx1514, A0=>nx1510, A1=>nx1517);
   ix107 : nor02ii port map ( Y=>nx947, A0=>nx1533, A1=>clk_cnt_6);
   ix1531 : or04 port map ( Y=>nx1530, A0=>nx1711, A1=>nx1701, A2=>nx947, A3
      =>nx1705);
   ix93 : nor02ii port map ( Y=>nx1711, A0=>clk_cnt_6, A1=>nx1533);
   ix75 : nor02ii port map ( Y=>nx943, A0=>nx1549, A1=>clk_cnt_4);
   ix1547 : or04 port map ( Y=>nx1546, A0=>nx1713, A1=>nx1701, A2=>nx943, A3
      =>nx1705);
   ix61 : nor02ii port map ( Y=>nx1713, A0=>clk_cnt_4, A1=>nx1549);
   ix1002 : mux21 port map ( Y=>nx1001, A0=>clk_cnt_1, A1=>nx18, S0=>nx1721
   );
   ix19 : nor02ii port map ( Y=>nx18, A0=>nx1572, A1=>nx0);
   ix992 : mux21 port map ( Y=>nx991, A0=>clk_cnt_0, A1=>nx4, S0=>nx1721);
   ix5 : nor02ii port map ( Y=>nx4, A0=>clk_cnt_0, A1=>nx0);
   ix1578 : or02 port map ( Y=>nx937, A0=>nx1699, A1=>nx610);
   ix515 : and03 port map ( Y=>nx514, A0=>nx1374, A1=>nx1357, A2=>nx1368);
   ix527 : and03 port map ( Y=>nx526, A0=>nx1402, A1=>nx1385, A2=>nx1391);
   ix537 : and03 port map ( Y=>nx536, A0=>nx1425, A1=>nx1408, A2=>nx1419);
   ix551 : and03 port map ( Y=>nx550, A0=>nx1453, A1=>nx1436, A2=>nx1442);
   ix561 : and03 port map ( Y=>nx560, A0=>nx1476, A1=>nx1459, A2=>nx1470);
   ix573 : and03 port map ( Y=>nx572, A0=>nx1504, A1=>nx1487, A2=>nx1493);
   ix583 : ao21 port map ( Y=>nx582, A0=>nx1562, A1=>nx1567, B0=>nx1553);
   ix589 : and02 port map ( Y=>nx588, A0=>nx1537, A1=>nx1543);
   ix1300 : and03 port map ( Y=>nx1299, A0=>nx0, A1=>nx1715, A2=>nx1721);
   ix1612 : xnor2 port map ( Y=>nx1715, A0=>nx1608, A1=>nx478);
   ix479 : nor02ii port map ( Y=>nx478, A0=>nx1327, A1=>clk_cnt_30);
   ix1616 : nor02ii port map ( Y=>nx1615, A0=>nx652, A1=>nx1608);
   ix653 : and04 port map ( Y=>nx652, A0=>nx1543, A1=>nx1527, A2=>nx1537, A3
      =>nx1717);
   ix1619 : and03 port map ( Y=>nx1717, A0=>nx644, A1=>nx1553, A2=>nx610);
   ix1718 : inv01 port map ( Y=>nx1719, A=>nx1705);
   ix1720 : inv01 port map ( Y=>nx1721, A=>nx1705);
end structural ;

