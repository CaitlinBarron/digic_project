//
// Verilog description for cell MAC, 
// Sun Dec  8 19:33:49 2019
//
// LeonardoSpectrum Level 3, 2008b.3 
//


module MAC ( A, B, clk, rst, test_mode, Result_OUT ) ;

    input [15:0]A ;
    input [15:0]B ;
    input clk ;
    input rst ;
    input test_mode ;
    output [31:0]Result_OUT ;

    wire MultIn1_15, MultIn1_14, MultIn1_13, MultIn1_12, MultIn1_11, MultIn1_10, 
         MultIn1_9, MultIn1_8, MultIn1_7, MultIn1_6, MultIn1_5, MultIn1_4, 
         MultIn1_3, MultIn1_2, MultIn1_1, MultIn1_0, MultIn2_15, MultIn2_14, 
         MultIn2_13, MultIn2_12, MultIn2_11, MultIn2_10, MultIn2_9, MultIn2_8, 
         MultIn2_7, MultIn2_6, MultIn2_5, MultIn2_4, MultIn2_3, MultIn2_2, 
         MultIn2_1, MultIn2_0, LFSR_OUT_31, LFSR_OUT_30, LFSR_OUT_29, 
         LFSR_OUT_28, LFSR_OUT_27, LFSR_OUT_26, LFSR_OUT_25, LFSR_OUT_24, 
         LFSR_OUT_23, LFSR_OUT_22, LFSR_OUT_21, LFSR_OUT_20, LFSR_OUT_19, 
         LFSR_OUT_18, LFSR_OUT_17, LFSR_OUT_16, LFSR_OUT_15, LFSR_OUT_14, 
         LFSR_OUT_13, LFSR_OUT_12, LFSR_OUT_11, LFSR_OUT_10, LFSR_OUT_9, 
         LFSR_OUT_8, LFSR_OUT_7, LFSR_OUT_6, LFSR_OUT_5, LFSR_OUT_4, LFSR_OUT_3, 
         LFSR_OUT_2, LFSR_OUT_1, LFSR_OUT_0, MISR_OUT_31, MISR_OUT_30, 
         MISR_OUT_29, MISR_OUT_28, MISR_OUT_27, MISR_OUT_26, MISR_OUT_25, 
         MISR_OUT_24, MISR_OUT_23, MISR_OUT_22, MISR_OUT_21, MISR_OUT_20, 
         MISR_OUT_19, MISR_OUT_18, MISR_OUT_17, MISR_OUT_16, MISR_OUT_15, 
         MISR_OUT_14, MISR_OUT_13, MISR_OUT_12, MISR_OUT_11, MISR_OUT_10, 
         MISR_OUT_9, MISR_OUT_8, MISR_OUT_7, MISR_OUT_6, MISR_OUT_5, MISR_OUT_4, 
         MISR_OUT_3, MISR_OUT_2, MISR_OUT_1, MISR_OUT_0, MULT_OUT_31, 
         MULT_OUT_30, MULT_OUT_29, MULT_OUT_28, MULT_OUT_27, MULT_OUT_26, 
         MULT_OUT_25, MULT_OUT_24, MULT_OUT_23, MULT_OUT_22, MULT_OUT_21, 
         MULT_OUT_20, MULT_OUT_19, MULT_OUT_18, MULT_OUT_17, MULT_OUT_16, 
         MULT_OUT_15, MULT_OUT_14, MULT_OUT_13, MULT_OUT_12, MULT_OUT_11, 
         MULT_OUT_10, MULT_OUT_9, MULT_OUT_8, MULT_OUT_7, MULT_OUT_6, MULT_OUT_5, 
         MULT_OUT_4, MULT_OUT_3, MULT_OUT_2, MULT_OUT_1, MULT_OUT_0, 
         ADDER_OUT_31, ADDER_OUT_30, ADDER_OUT_29, ADDER_OUT_28, ADDER_OUT_27, 
         ADDER_OUT_26, ADDER_OUT_25, ADDER_OUT_24, ADDER_OUT_23, ADDER_OUT_22, 
         ADDER_OUT_21, ADDER_OUT_20, ADDER_OUT_19, ADDER_OUT_18, ADDER_OUT_17, 
         ADDER_OUT_16, ADDER_OUT_15, ADDER_OUT_14, ADDER_OUT_13, ADDER_OUT_12, 
         ADDER_OUT_11, ADDER_OUT_10, ADDER_OUT_9, ADDER_OUT_8, ADDER_OUT_7, 
         ADDER_OUT_6, ADDER_OUT_5, ADDER_OUT_4, ADDER_OUT_3, ADDER_OUT_2, 
         ADDER_OUT_1, ADDER_OUT_0, REG_OUT_31, REG_OUT_30, REG_OUT_29, 
         REG_OUT_28, REG_OUT_27, REG_OUT_26, REG_OUT_25, REG_OUT_24, REG_OUT_23, 
         REG_OUT_22, REG_OUT_21, REG_OUT_20, REG_OUT_19, REG_OUT_18, REG_OUT_17, 
         REG_OUT_16, REG_OUT_15, REG_OUT_14, REG_OUT_13, REG_OUT_12, REG_OUT_11, 
         REG_OUT_10, REG_OUT_9, REG_OUT_8, REG_OUT_7, REG_OUT_6, REG_OUT_5, 
         REG_OUT_4, REG_OUT_3, REG_OUT_2, REG_OUT_1, REG_OUT_0, MISR_EN, GND0, 
         PWR, nx0, clk_cnt_30, nx937, clk_cnt_29, clk_cnt_28, clk_cnt_27, 
         clk_cnt_26, clk_cnt_25, clk_cnt_24, clk_cnt_23, clk_cnt_22, clk_cnt_21, 
         clk_cnt_20, clk_cnt_19, clk_cnt_18, clk_cnt_17, clk_cnt_16, clk_cnt_15, 
         clk_cnt_14, clk_cnt_13, clk_cnt_12, clk_cnt_11, clk_cnt_10, clk_cnt_9, 
         clk_cnt_8, clk_cnt_7, clk_cnt_6, clk_cnt_5, clk_cnt_4, clk_cnt_3, 
         clk_cnt_2, clk_cnt_1, clk_cnt_0, nx4, nx18, nx28, nx44, nx943, nx76, 
         nx947, nx108, nx949, nx130, nx140, nx953, nx162, nx172, nx956, nx194, 
         nx204, nx959, nx226, nx236, nx963, nx258, nx268, nx965, nx290, nx300, 
         nx969, nx322, nx332, nx972, nx354, nx364, nx975, nx386, nx396, nx979, 
         nx418, nx428, nx981, nx450, nx460, nx478, nx484, nx504, nx514, nx526, 
         nx536, nx550, nx560, nx572, nx582, nx588, nx602, nx610, nx644, nx652, 
         nx662, nx991, nx1001, nx1011, nx1021, nx1031, nx1041, nx1051, nx1061, 
         nx1071, nx1081, nx1091, nx1101, nx1111, nx1121, nx1131, nx1141, nx1151, 
         nx1161, nx1171, nx1181, nx1191, nx1201, nx1211, nx1221, nx1231, nx1241, 
         nx1251, nx1261, nx1271, nx1281, nx1291, nx1299, nx1311, nx1321, nx1327, 
         nx1331, nx1334, nx1336, nx1340, nx1344, nx1347, nx1351, nx1353, nx1357, 
         nx1361, nx1364, nx1368, nx1370, nx1374, nx1378, nx1381, nx1385, nx1387, 
         nx1391, nx1395, nx1398, nx1402, nx1404, nx1408, nx1412, nx1415, nx1419, 
         nx1421, nx1425, nx1429, nx1432, nx1436, nx1438, nx1442, nx1446, nx1449, 
         nx1453, nx1455, nx1459, nx1463, nx1466, nx1470, nx1472, nx1476, nx1480, 
         nx1483, nx1487, nx1489, nx1493, nx1497, nx1500, nx1504, nx1506, nx1510, 
         nx1514, nx1517, nx1521, nx1523, nx1527, nx1530, nx1533, nx1537, nx1539, 
         nx1543, nx1546, nx1549, nx1553, nx1555, nx1558, nx1562, nx1564, nx1567, 
         nx1572, nx1590, nx1592, nx1597, nx1603, nx1608, nx1615, nx1691, nx1693, 
         nx1695, nx1697, nx1699, nx1701, nx1705, nx1711, nx1713, nx1715, nx1717, 
         nx1719, nx1721;
    wire [4:0] \$dummy ;




    Multiplier_32 Multiplier0 (.A ({MultIn1_15,MultIn1_14,MultIn1_13,MultIn1_12,
                  MultIn1_11,MultIn1_10,MultIn1_9,MultIn1_8,MultIn1_7,MultIn1_6,
                  MultIn1_5,MultIn1_4,MultIn1_3,MultIn1_2,MultIn1_1,MultIn1_0})
                  , .B ({MultIn2_15,MultIn2_14,MultIn2_13,MultIn2_12,MultIn2_11,
                  MultIn2_10,MultIn2_9,MultIn2_8,MultIn2_7,MultIn2_6,MultIn2_5,
                  MultIn2_4,MultIn2_3,MultIn2_2,MultIn2_1,MultIn2_0}), .Product (
                  {MULT_OUT_31,MULT_OUT_30,MULT_OUT_29,MULT_OUT_28,MULT_OUT_27,
                  MULT_OUT_26,MULT_OUT_25,MULT_OUT_24,MULT_OUT_23,MULT_OUT_22,
                  MULT_OUT_21,MULT_OUT_20,MULT_OUT_19,MULT_OUT_18,MULT_OUT_17,
                  MULT_OUT_16,MULT_OUT_15,MULT_OUT_14,MULT_OUT_13,MULT_OUT_12,
                  MULT_OUT_11,MULT_OUT_10,MULT_OUT_9,MULT_OUT_8,MULT_OUT_7,
                  MULT_OUT_6,MULT_OUT_5,MULT_OUT_4,MULT_OUT_3,MULT_OUT_2,
                  MULT_OUT_1,MULT_OUT_0})) ;
    RegisterN_32 RegisterN0 (.clk (clk), .reset (rst), .enable (PWR), .\input  (
                 {ADDER_OUT_31,ADDER_OUT_30,ADDER_OUT_29,ADDER_OUT_28,
                 ADDER_OUT_27,ADDER_OUT_26,ADDER_OUT_25,ADDER_OUT_24,
                 ADDER_OUT_23,ADDER_OUT_22,ADDER_OUT_21,ADDER_OUT_20,
                 ADDER_OUT_19,ADDER_OUT_18,ADDER_OUT_17,ADDER_OUT_16,
                 ADDER_OUT_15,ADDER_OUT_14,ADDER_OUT_13,ADDER_OUT_12,
                 ADDER_OUT_11,ADDER_OUT_10,ADDER_OUT_9,ADDER_OUT_8,ADDER_OUT_7,
                 ADDER_OUT_6,ADDER_OUT_5,ADDER_OUT_4,ADDER_OUT_3,ADDER_OUT_2,
                 ADDER_OUT_1,ADDER_OUT_0}), .\output  ({REG_OUT_31,REG_OUT_30,
                 REG_OUT_29,REG_OUT_28,REG_OUT_27,REG_OUT_26,REG_OUT_25,
                 REG_OUT_24,REG_OUT_23,REG_OUT_22,REG_OUT_21,REG_OUT_20,
                 REG_OUT_19,REG_OUT_18,REG_OUT_17,REG_OUT_16,REG_OUT_15,
                 REG_OUT_14,REG_OUT_13,REG_OUT_12,REG_OUT_11,REG_OUT_10,
                 REG_OUT_9,REG_OUT_8,REG_OUT_7,REG_OUT_6,REG_OUT_5,REG_OUT_4,
                 REG_OUT_3,REG_OUT_2,REG_OUT_1,REG_OUT_0})) ;
    LFSR LFSR0 (.clk (clk), .rst (rst), .enable (test_mode), .bit_pattern ({
         LFSR_OUT_31,LFSR_OUT_30,LFSR_OUT_29,LFSR_OUT_28,LFSR_OUT_27,LFSR_OUT_26
         ,LFSR_OUT_25,LFSR_OUT_24,LFSR_OUT_23,LFSR_OUT_22,LFSR_OUT_21,
         LFSR_OUT_20,LFSR_OUT_19,LFSR_OUT_18,LFSR_OUT_17,LFSR_OUT_16,LFSR_OUT_15
         ,LFSR_OUT_14,LFSR_OUT_13,LFSR_OUT_12,LFSR_OUT_11,LFSR_OUT_10,LFSR_OUT_9
         ,LFSR_OUT_8,LFSR_OUT_7,LFSR_OUT_6,LFSR_OUT_5,LFSR_OUT_4,LFSR_OUT_3,
         LFSR_OUT_2,LFSR_OUT_1,LFSR_OUT_0})) ;
    MISR MISR0 (.clk (clk), .rst (rst), .enable (MISR_EN), .mult_result ({
         REG_OUT_31,REG_OUT_30,REG_OUT_29,REG_OUT_28,REG_OUT_27,REG_OUT_26,
         REG_OUT_25,REG_OUT_24,REG_OUT_23,REG_OUT_22,REG_OUT_21,REG_OUT_20,
         REG_OUT_19,REG_OUT_18,REG_OUT_17,REG_OUT_16,REG_OUT_15,REG_OUT_14,
         REG_OUT_13,REG_OUT_12,REG_OUT_11,REG_OUT_10,REG_OUT_9,REG_OUT_8,
         REG_OUT_7,REG_OUT_6,REG_OUT_5,REG_OUT_4,REG_OUT_3,REG_OUT_2,REG_OUT_1,
         REG_OUT_0}), .signature ({MISR_OUT_31,MISR_OUT_30,MISR_OUT_29,
         MISR_OUT_28,MISR_OUT_27,MISR_OUT_26,MISR_OUT_25,MISR_OUT_24,MISR_OUT_23
         ,MISR_OUT_22,MISR_OUT_21,MISR_OUT_20,MISR_OUT_19,MISR_OUT_18,
         MISR_OUT_17,MISR_OUT_16,MISR_OUT_15,MISR_OUT_14,MISR_OUT_13,MISR_OUT_12
         ,MISR_OUT_11,MISR_OUT_10,MISR_OUT_9,MISR_OUT_8,MISR_OUT_7,MISR_OUT_6,
         MISR_OUT_5,MISR_OUT_4,MISR_OUT_3,MISR_OUT_2,MISR_OUT_1,MISR_OUT_0})) ;
    RCFA_32 RCFA0 (.A ({MULT_OUT_31,MULT_OUT_30,MULT_OUT_29,MULT_OUT_28,
            MULT_OUT_27,MULT_OUT_26,MULT_OUT_25,MULT_OUT_24,MULT_OUT_23,
            MULT_OUT_22,MULT_OUT_21,MULT_OUT_20,MULT_OUT_19,MULT_OUT_18,
            MULT_OUT_17,MULT_OUT_16,MULT_OUT_15,MULT_OUT_14,MULT_OUT_13,
            MULT_OUT_12,MULT_OUT_11,MULT_OUT_10,MULT_OUT_9,MULT_OUT_8,MULT_OUT_7
            ,MULT_OUT_6,MULT_OUT_5,MULT_OUT_4,MULT_OUT_3,MULT_OUT_2,MULT_OUT_1,
            MULT_OUT_0}), .B ({REG_OUT_31,REG_OUT_30,REG_OUT_29,REG_OUT_28,
            REG_OUT_27,REG_OUT_26,REG_OUT_25,REG_OUT_24,REG_OUT_23,REG_OUT_22,
            REG_OUT_21,REG_OUT_20,REG_OUT_19,REG_OUT_18,REG_OUT_17,REG_OUT_16,
            REG_OUT_15,REG_OUT_14,REG_OUT_13,REG_OUT_12,REG_OUT_11,REG_OUT_10,
            REG_OUT_9,REG_OUT_8,REG_OUT_7,REG_OUT_6,REG_OUT_5,REG_OUT_4,
            REG_OUT_3,REG_OUT_2,REG_OUT_1,REG_OUT_0}), .Cin (GND0), .Sum ({
            ADDER_OUT_31,ADDER_OUT_30,ADDER_OUT_29,ADDER_OUT_28,ADDER_OUT_27,
            ADDER_OUT_26,ADDER_OUT_25,ADDER_OUT_24,ADDER_OUT_23,ADDER_OUT_22,
            ADDER_OUT_21,ADDER_OUT_20,ADDER_OUT_19,ADDER_OUT_18,ADDER_OUT_17,
            ADDER_OUT_16,ADDER_OUT_15,ADDER_OUT_14,ADDER_OUT_13,ADDER_OUT_12,
            ADDER_OUT_11,ADDER_OUT_10,ADDER_OUT_9,ADDER_OUT_8,ADDER_OUT_7,
            ADDER_OUT_6,ADDER_OUT_5,ADDER_OUT_4,ADDER_OUT_3,ADDER_OUT_2,
            ADDER_OUT_1,ADDER_OUT_0}), .Cout (\$dummy [0])) ;
    fake_vcc ix799 (.Y (PWR)) ;
    fake_gnd ix797 (.Y (GND0)) ;
    dff reg_MISR_EN (.Q (MISR_EN), .QB (\$dummy [1]), .D (nx1311), .CLK (clk)) ;
    mux21 ix663 (.Y (nx662), .A0 (MISR_EN), .A1 (nx610), .S0 (nx1615)) ;
    oai21 ix611 (.Y (nx610), .A0 (nx1321), .A1 (nx1597), .B0 (nx1608)) ;
    nand04 ix1322 (.Y (nx1321), .A0 (nx504), .A1 (nx514), .A2 (nx526), .A3 (
           nx536)) ;
    aoi21 ix485 (.Y (nx484), .A0 (nx1327), .A1 (nx1590), .B0 (nx1592)) ;
    nand02 ix1328 (.Y (nx1327), .A0 (clk_cnt_29), .A1 (nx981)) ;
    oai21 ix1282 (.Y (nx1281), .A0 (nx1331), .A1 (nx1693), .B0 (nx1336)) ;
    dff reg_clk_cnt_29 (.Q (clk_cnt_29), .QB (nx1331), .D (nx1281), .CLK (clk)
        ) ;
    nand02 ix1335 (.Y (nx1334), .A0 (rst), .A1 (test_mode)) ;
    nand04 ix1337 (.Y (nx1336), .A0 (nx460), .A1 (nx0), .A2 (nx1327), .A3 (
           nx1697)) ;
    or02 ix461 (.Y (nx460), .A0 (nx981), .A1 (clk_cnt_29)) ;
    nor03 ix451 (.Y (nx450), .A0 (nx1344), .A1 (nx1699), .A2 (nx981)) ;
    dff reg_clk_cnt_28 (.Q (clk_cnt_28), .QB (nx1340), .D (nx1271), .CLK (clk)
        ) ;
    nand02 ix1348 (.Y (nx1347), .A0 (clk_cnt_27), .A1 (nx979)) ;
    oai21 ix1262 (.Y (nx1261), .A0 (nx1351), .A1 (nx1693), .B0 (nx1353)) ;
    dff reg_clk_cnt_27 (.Q (clk_cnt_27), .QB (nx1351), .D (nx1261), .CLK (clk)
        ) ;
    nand04 ix1354 (.Y (nx1353), .A0 (nx428), .A1 (nx0), .A2 (nx1347), .A3 (
           nx1697)) ;
    or02 ix429 (.Y (nx428), .A0 (nx979), .A1 (clk_cnt_27)) ;
    nor03 ix419 (.Y (nx418), .A0 (nx1361), .A1 (nx1699), .A2 (nx979)) ;
    dff reg_clk_cnt_26 (.Q (clk_cnt_26), .QB (nx1357), .D (nx1251), .CLK (clk)
        ) ;
    nand02 ix1365 (.Y (nx1364), .A0 (clk_cnt_25), .A1 (nx975)) ;
    oai21 ix1242 (.Y (nx1241), .A0 (nx1368), .A1 (nx1693), .B0 (nx1370)) ;
    dff reg_clk_cnt_25 (.Q (clk_cnt_25), .QB (nx1368), .D (nx1241), .CLK (clk)
        ) ;
    nand04 ix1371 (.Y (nx1370), .A0 (nx396), .A1 (nx0), .A2 (nx1364), .A3 (
           nx1697)) ;
    or02 ix397 (.Y (nx396), .A0 (nx975), .A1 (clk_cnt_25)) ;
    nor03 ix387 (.Y (nx386), .A0 (nx1378), .A1 (nx1699), .A2 (nx975)) ;
    dff reg_clk_cnt_24 (.Q (clk_cnt_24), .QB (nx1374), .D (nx1231), .CLK (clk)
        ) ;
    nand02 ix1382 (.Y (nx1381), .A0 (clk_cnt_23), .A1 (nx972)) ;
    oai21 ix1222 (.Y (nx1221), .A0 (nx1385), .A1 (nx1693), .B0 (nx1387)) ;
    dff reg_clk_cnt_23 (.Q (clk_cnt_23), .QB (nx1385), .D (nx1221), .CLK (clk)
        ) ;
    nand04 ix1388 (.Y (nx1387), .A0 (nx364), .A1 (nx0), .A2 (nx1381), .A3 (
           nx1697)) ;
    or02 ix365 (.Y (nx364), .A0 (nx972), .A1 (clk_cnt_23)) ;
    nor03 ix355 (.Y (nx354), .A0 (nx1395), .A1 (nx1699), .A2 (nx972)) ;
    dff reg_clk_cnt_22 (.Q (clk_cnt_22), .QB (nx1391), .D (nx1211), .CLK (clk)
        ) ;
    nand02 ix1399 (.Y (nx1398), .A0 (clk_cnt_21), .A1 (nx969)) ;
    oai21 ix1202 (.Y (nx1201), .A0 (nx1402), .A1 (nx1693), .B0 (nx1404)) ;
    dff reg_clk_cnt_21 (.Q (clk_cnt_21), .QB (nx1402), .D (nx1201), .CLK (clk)
        ) ;
    nand04 ix1405 (.Y (nx1404), .A0 (nx332), .A1 (nx1691), .A2 (nx1398), .A3 (
           nx1695)) ;
    or02 ix333 (.Y (nx332), .A0 (nx969), .A1 (clk_cnt_21)) ;
    nor03 ix323 (.Y (nx322), .A0 (nx1412), .A1 (nx1699), .A2 (nx969)) ;
    dff reg_clk_cnt_20 (.Q (clk_cnt_20), .QB (nx1408), .D (nx1191), .CLK (clk)
        ) ;
    nand02 ix1416 (.Y (nx1415), .A0 (clk_cnt_19), .A1 (nx965)) ;
    oai21 ix1182 (.Y (nx1181), .A0 (nx1419), .A1 (nx1693), .B0 (nx1421)) ;
    dff reg_clk_cnt_19 (.Q (clk_cnt_19), .QB (nx1419), .D (nx1181), .CLK (clk)
        ) ;
    nand04 ix1422 (.Y (nx1421), .A0 (nx300), .A1 (nx1691), .A2 (nx1415), .A3 (
           nx1695)) ;
    or02 ix301 (.Y (nx300), .A0 (nx965), .A1 (clk_cnt_19)) ;
    nor03 ix291 (.Y (nx290), .A0 (nx1429), .A1 (nx1699), .A2 (nx965)) ;
    dff reg_clk_cnt_18 (.Q (clk_cnt_18), .QB (nx1425), .D (nx1171), .CLK (clk)
        ) ;
    nand02 ix1433 (.Y (nx1432), .A0 (clk_cnt_17), .A1 (nx963)) ;
    oai21 ix1162 (.Y (nx1161), .A0 (nx1436), .A1 (nx1693), .B0 (nx1438)) ;
    dff reg_clk_cnt_17 (.Q (clk_cnt_17), .QB (nx1436), .D (nx1161), .CLK (clk)
        ) ;
    nand04 ix1439 (.Y (nx1438), .A0 (nx268), .A1 (nx1691), .A2 (nx1432), .A3 (
           nx1695)) ;
    or02 ix269 (.Y (nx268), .A0 (nx963), .A1 (clk_cnt_17)) ;
    nor03 ix259 (.Y (nx258), .A0 (nx1446), .A1 (nx1699), .A2 (nx963)) ;
    dff reg_clk_cnt_16 (.Q (clk_cnt_16), .QB (nx1442), .D (nx1151), .CLK (clk)
        ) ;
    nand02 ix1450 (.Y (nx1449), .A0 (clk_cnt_15), .A1 (nx959)) ;
    oai21 ix1142 (.Y (nx1141), .A0 (nx1453), .A1 (nx1693), .B0 (nx1455)) ;
    dff reg_clk_cnt_15 (.Q (clk_cnt_15), .QB (nx1453), .D (nx1141), .CLK (clk)
        ) ;
    nand04 ix1456 (.Y (nx1455), .A0 (nx236), .A1 (nx1691), .A2 (nx1449), .A3 (
           nx1695)) ;
    or02 ix237 (.Y (nx236), .A0 (nx959), .A1 (clk_cnt_15)) ;
    nor03 ix227 (.Y (nx226), .A0 (nx1463), .A1 (nx1699), .A2 (nx959)) ;
    dff reg_clk_cnt_14 (.Q (clk_cnt_14), .QB (nx1459), .D (nx1131), .CLK (clk)
        ) ;
    nand02 ix1467 (.Y (nx1466), .A0 (clk_cnt_13), .A1 (nx956)) ;
    oai21 ix1122 (.Y (nx1121), .A0 (nx1470), .A1 (nx1693), .B0 (nx1472)) ;
    dff reg_clk_cnt_13 (.Q (clk_cnt_13), .QB (nx1470), .D (nx1121), .CLK (clk)
        ) ;
    nand04 ix1473 (.Y (nx1472), .A0 (nx204), .A1 (nx1691), .A2 (nx1466), .A3 (
           nx1695)) ;
    or02 ix205 (.Y (nx204), .A0 (nx956), .A1 (clk_cnt_13)) ;
    nor03 ix195 (.Y (nx194), .A0 (nx1480), .A1 (nx1699), .A2 (nx956)) ;
    dff reg_clk_cnt_12 (.Q (clk_cnt_12), .QB (nx1476), .D (nx1111), .CLK (clk)
        ) ;
    nand02 ix1484 (.Y (nx1483), .A0 (clk_cnt_11), .A1 (nx953)) ;
    oai21 ix1102 (.Y (nx1101), .A0 (nx1487), .A1 (nx1693), .B0 (nx1489)) ;
    dff reg_clk_cnt_11 (.Q (clk_cnt_11), .QB (nx1487), .D (nx1101), .CLK (clk)
        ) ;
    nand04 ix1490 (.Y (nx1489), .A0 (nx172), .A1 (nx1691), .A2 (nx1483), .A3 (
           nx1695)) ;
    or02 ix173 (.Y (nx172), .A0 (nx953), .A1 (clk_cnt_11)) ;
    nor03 ix163 (.Y (nx162), .A0 (nx1497), .A1 (nx1699), .A2 (nx953)) ;
    dff reg_clk_cnt_10 (.Q (clk_cnt_10), .QB (nx1493), .D (nx1091), .CLK (clk)
        ) ;
    nand02 ix1501 (.Y (nx1500), .A0 (clk_cnt_9), .A1 (nx949)) ;
    oai21 ix1082 (.Y (nx1081), .A0 (nx1504), .A1 (nx1693), .B0 (nx1506)) ;
    dff reg_clk_cnt_9 (.Q (clk_cnt_9), .QB (nx1504), .D (nx1081), .CLK (clk)) ;
    nand04 ix1507 (.Y (nx1506), .A0 (nx140), .A1 (nx1691), .A2 (nx1500), .A3 (
           nx1695)) ;
    or02 ix141 (.Y (nx140), .A0 (nx949), .A1 (clk_cnt_9)) ;
    nor03 ix131 (.Y (nx130), .A0 (nx1514), .A1 (nx1699), .A2 (nx949)) ;
    dff reg_clk_cnt_8 (.Q (clk_cnt_8), .QB (nx1510), .D (nx1071), .CLK (clk)) ;
    nand02 ix1518 (.Y (nx1517), .A0 (clk_cnt_7), .A1 (nx947)) ;
    oai21 ix1062 (.Y (nx1061), .A0 (nx1521), .A1 (nx1693), .B0 (nx1523)) ;
    dff reg_clk_cnt_7 (.Q (clk_cnt_7), .QB (nx1521), .D (nx1061), .CLK (clk)) ;
    nand04 ix1524 (.Y (nx1523), .A0 (nx108), .A1 (nx1691), .A2 (nx1517), .A3 (
           nx1695)) ;
    or02 ix109 (.Y (nx108), .A0 (nx947), .A1 (clk_cnt_7)) ;
    oai21 ix1052 (.Y (nx1051), .A0 (nx1527), .A1 (nx1693), .B0 (nx1530)) ;
    nand02 ix1534 (.Y (nx1533), .A0 (clk_cnt_5), .A1 (nx943)) ;
    oai21 ix1042 (.Y (nx1041), .A0 (nx1537), .A1 (nx1693), .B0 (nx1539)) ;
    dff reg_clk_cnt_5 (.Q (clk_cnt_5), .QB (nx1537), .D (nx1041), .CLK (clk)) ;
    nand04 ix1540 (.Y (nx1539), .A0 (nx76), .A1 (nx1691), .A2 (nx1533), .A3 (
           nx1695)) ;
    or02 ix77 (.Y (nx76), .A0 (nx943), .A1 (clk_cnt_5)) ;
    oai21 ix1032 (.Y (nx1031), .A0 (nx1543), .A1 (nx1693), .B0 (nx1546)) ;
    nand04 ix1550 (.Y (nx1549), .A0 (clk_cnt_3), .A1 (clk_cnt_2), .A2 (clk_cnt_1
           ), .A3 (clk_cnt_0)) ;
    oai21 ix1022 (.Y (nx1021), .A0 (nx1553), .A1 (nx1695), .B0 (nx1555)) ;
    dff reg_clk_cnt_3 (.Q (clk_cnt_3), .QB (nx1553), .D (nx1021), .CLK (clk)) ;
    nand04 ix1556 (.Y (nx1555), .A0 (nx44), .A1 (nx1691), .A2 (nx1549), .A3 (
           nx1695)) ;
    nand02 ix45 (.Y (nx44), .A0 (nx1558), .A1 (nx1553)) ;
    nand03 ix1559 (.Y (nx1558), .A0 (clk_cnt_2), .A1 (clk_cnt_1), .A2 (clk_cnt_0
           )) ;
    oai21 ix1012 (.Y (nx1011), .A0 (nx1562), .A1 (nx1695), .B0 (nx1564)) ;
    dff reg_clk_cnt_2 (.Q (clk_cnt_2), .QB (nx1562), .D (nx1011), .CLK (clk)) ;
    nand04 ix1565 (.Y (nx1564), .A0 (nx28), .A1 (nx1691), .A2 (nx1558), .A3 (
           nx1695)) ;
    nand02 ix29 (.Y (nx28), .A0 (nx1567), .A1 (nx1562)) ;
    nand02 ix1568 (.Y (nx1567), .A0 (clk_cnt_1), .A1 (clk_cnt_0)) ;
    dff reg_clk_cnt_1 (.Q (clk_cnt_1), .QB (\$dummy [2]), .D (nx1001), .CLK (clk
        )) ;
    oai21 ix1573 (.Y (nx1572), .A0 (clk_cnt_0), .A1 (clk_cnt_1), .B0 (nx1567)) ;
    dff reg_clk_cnt_0 (.Q (clk_cnt_0), .QB (\$dummy [3]), .D (nx991), .CLK (clk)
        ) ;
    dff reg_clk_cnt_4 (.Q (clk_cnt_4), .QB (nx1543), .D (nx1031), .CLK (clk)) ;
    dff reg_clk_cnt_6 (.Q (clk_cnt_6), .QB (nx1527), .D (nx1051), .CLK (clk)) ;
    dff reg_clk_cnt_30 (.Q (clk_cnt_30), .QB (nx1590), .D (nx1291), .CLK (clk)
        ) ;
    oai21 ix1593 (.Y (nx1592), .A0 (nx1590), .A1 (nx1327), .B0 (nx1691)) ;
    nand04 ix1598 (.Y (nx1597), .A0 (nx550), .A1 (nx560), .A2 (nx572), .A3 (
           nx602)) ;
    nor03 ix603 (.Y (nx602), .A0 (nx1603), .A1 (clk_cnt_8), .A2 (clk_cnt_7)) ;
    aoi21 ix1604 (.Y (nx1603), .A0 (nx582), .A1 (nx588), .B0 (nx1527)) ;
    dff clk_cnt_31 (.Q (\$dummy [4]), .QB (nx1608), .D (nx1299), .CLK (clk)) ;
    oai21 ix645 (.Y (nx644), .A0 (clk_cnt_1), .A1 (clk_cnt_0), .B0 (clk_cnt_2)
          ) ;
    mux21 ix805 (.Y (MultIn2_0), .A0 (B[0]), .A1 (LFSR_OUT_0), .S0 (test_mode)
          ) ;
    mux21 ix813 (.Y (MultIn2_1), .A0 (B[1]), .A1 (LFSR_OUT_1), .S0 (test_mode)
          ) ;
    mux21 ix821 (.Y (MultIn2_2), .A0 (B[2]), .A1 (LFSR_OUT_2), .S0 (test_mode)
          ) ;
    mux21 ix829 (.Y (MultIn2_3), .A0 (B[3]), .A1 (LFSR_OUT_3), .S0 (test_mode)
          ) ;
    mux21 ix837 (.Y (MultIn2_4), .A0 (B[4]), .A1 (LFSR_OUT_4), .S0 (test_mode)
          ) ;
    mux21 ix845 (.Y (MultIn2_5), .A0 (B[5]), .A1 (LFSR_OUT_5), .S0 (test_mode)
          ) ;
    mux21 ix853 (.Y (MultIn2_6), .A0 (B[6]), .A1 (LFSR_OUT_6), .S0 (test_mode)
          ) ;
    mux21 ix861 (.Y (MultIn2_7), .A0 (B[7]), .A1 (LFSR_OUT_7), .S0 (test_mode)
          ) ;
    mux21 ix869 (.Y (MultIn2_8), .A0 (B[8]), .A1 (LFSR_OUT_8), .S0 (test_mode)
          ) ;
    mux21 ix877 (.Y (MultIn2_9), .A0 (B[9]), .A1 (LFSR_OUT_9), .S0 (test_mode)
          ) ;
    mux21 ix885 (.Y (MultIn2_10), .A0 (B[10]), .A1 (LFSR_OUT_10), .S0 (test_mode
          )) ;
    mux21 ix893 (.Y (MultIn2_11), .A0 (B[11]), .A1 (LFSR_OUT_11), .S0 (test_mode
          )) ;
    mux21 ix901 (.Y (MultIn2_12), .A0 (B[12]), .A1 (LFSR_OUT_12), .S0 (test_mode
          )) ;
    mux21 ix909 (.Y (MultIn2_13), .A0 (B[13]), .A1 (LFSR_OUT_13), .S0 (test_mode
          )) ;
    mux21 ix917 (.Y (MultIn2_14), .A0 (B[14]), .A1 (LFSR_OUT_14), .S0 (test_mode
          )) ;
    mux21 ix925 (.Y (MultIn2_15), .A0 (B[15]), .A1 (LFSR_OUT_15), .S0 (test_mode
          )) ;
    mux21 ix677 (.Y (MultIn1_0), .A0 (A[0]), .A1 (LFSR_OUT_16), .S0 (test_mode)
          ) ;
    mux21 ix685 (.Y (MultIn1_1), .A0 (A[1]), .A1 (LFSR_OUT_17), .S0 (test_mode)
          ) ;
    mux21 ix693 (.Y (MultIn1_2), .A0 (A[2]), .A1 (LFSR_OUT_18), .S0 (test_mode)
          ) ;
    mux21 ix701 (.Y (MultIn1_3), .A0 (A[3]), .A1 (LFSR_OUT_19), .S0 (test_mode)
          ) ;
    mux21 ix709 (.Y (MultIn1_4), .A0 (A[4]), .A1 (LFSR_OUT_20), .S0 (test_mode)
          ) ;
    mux21 ix717 (.Y (MultIn1_5), .A0 (A[5]), .A1 (LFSR_OUT_21), .S0 (test_mode)
          ) ;
    mux21 ix725 (.Y (MultIn1_6), .A0 (A[6]), .A1 (LFSR_OUT_22), .S0 (test_mode)
          ) ;
    mux21 ix733 (.Y (MultIn1_7), .A0 (A[7]), .A1 (LFSR_OUT_23), .S0 (test_mode)
          ) ;
    mux21 ix741 (.Y (MultIn1_8), .A0 (A[8]), .A1 (LFSR_OUT_24), .S0 (test_mode)
          ) ;
    mux21 ix749 (.Y (MultIn1_9), .A0 (A[9]), .A1 (LFSR_OUT_25), .S0 (test_mode)
          ) ;
    mux21 ix757 (.Y (MultIn1_10), .A0 (A[10]), .A1 (LFSR_OUT_26), .S0 (test_mode
          )) ;
    mux21 ix765 (.Y (MultIn1_11), .A0 (A[11]), .A1 (LFSR_OUT_27), .S0 (test_mode
          )) ;
    mux21 ix773 (.Y (MultIn1_12), .A0 (A[12]), .A1 (LFSR_OUT_28), .S0 (test_mode
          )) ;
    mux21 ix781 (.Y (MultIn1_13), .A0 (A[13]), .A1 (LFSR_OUT_29), .S0 (test_mode
          )) ;
    mux21 ix789 (.Y (MultIn1_14), .A0 (A[14]), .A1 (LFSR_OUT_30), .S0 (test_mode
          )) ;
    mux21 ix801 (.Y (MultIn1_15), .A0 (A[15]), .A1 (LFSR_OUT_31), .S0 (test_mode
          )) ;
    mux21 ix933 (.Y (Result_OUT[0]), .A0 (REG_OUT_0), .A1 (MISR_OUT_0), .S0 (
          test_mode)) ;
    mux21 ix941 (.Y (Result_OUT[1]), .A0 (REG_OUT_1), .A1 (MISR_OUT_1), .S0 (
          test_mode)) ;
    mux21 ix949 (.Y (Result_OUT[2]), .A0 (REG_OUT_2), .A1 (MISR_OUT_2), .S0 (
          test_mode)) ;
    mux21 ix957 (.Y (Result_OUT[3]), .A0 (REG_OUT_3), .A1 (MISR_OUT_3), .S0 (
          test_mode)) ;
    mux21 ix965 (.Y (Result_OUT[4]), .A0 (REG_OUT_4), .A1 (MISR_OUT_4), .S0 (
          test_mode)) ;
    mux21 ix973 (.Y (Result_OUT[5]), .A0 (REG_OUT_5), .A1 (MISR_OUT_5), .S0 (
          test_mode)) ;
    mux21 ix981 (.Y (Result_OUT[6]), .A0 (REG_OUT_6), .A1 (MISR_OUT_6), .S0 (
          test_mode)) ;
    mux21 ix989 (.Y (Result_OUT[7]), .A0 (REG_OUT_7), .A1 (MISR_OUT_7), .S0 (
          test_mode)) ;
    mux21 ix997 (.Y (Result_OUT[8]), .A0 (REG_OUT_8), .A1 (MISR_OUT_8), .S0 (
          test_mode)) ;
    mux21 ix1005 (.Y (Result_OUT[9]), .A0 (REG_OUT_9), .A1 (MISR_OUT_9), .S0 (
          test_mode)) ;
    mux21 ix1013 (.Y (Result_OUT[10]), .A0 (REG_OUT_10), .A1 (MISR_OUT_10), .S0 (
          test_mode)) ;
    mux21 ix1021 (.Y (Result_OUT[11]), .A0 (REG_OUT_11), .A1 (MISR_OUT_11), .S0 (
          test_mode)) ;
    mux21 ix1029 (.Y (Result_OUT[12]), .A0 (REG_OUT_12), .A1 (MISR_OUT_12), .S0 (
          test_mode)) ;
    mux21 ix1037 (.Y (Result_OUT[13]), .A0 (REG_OUT_13), .A1 (MISR_OUT_13), .S0 (
          test_mode)) ;
    mux21 ix1045 (.Y (Result_OUT[14]), .A0 (REG_OUT_14), .A1 (MISR_OUT_14), .S0 (
          test_mode)) ;
    mux21 ix1053 (.Y (Result_OUT[15]), .A0 (REG_OUT_15), .A1 (MISR_OUT_15), .S0 (
          test_mode)) ;
    mux21 ix1061 (.Y (Result_OUT[16]), .A0 (REG_OUT_16), .A1 (MISR_OUT_16), .S0 (
          test_mode)) ;
    mux21 ix1069 (.Y (Result_OUT[17]), .A0 (REG_OUT_17), .A1 (MISR_OUT_17), .S0 (
          test_mode)) ;
    mux21 ix1077 (.Y (Result_OUT[18]), .A0 (REG_OUT_18), .A1 (MISR_OUT_18), .S0 (
          test_mode)) ;
    mux21 ix1085 (.Y (Result_OUT[19]), .A0 (REG_OUT_19), .A1 (MISR_OUT_19), .S0 (
          test_mode)) ;
    mux21 ix1093 (.Y (Result_OUT[20]), .A0 (REG_OUT_20), .A1 (MISR_OUT_20), .S0 (
          test_mode)) ;
    mux21 ix1101 (.Y (Result_OUT[21]), .A0 (REG_OUT_21), .A1 (MISR_OUT_21), .S0 (
          test_mode)) ;
    mux21 ix1109 (.Y (Result_OUT[22]), .A0 (REG_OUT_22), .A1 (MISR_OUT_22), .S0 (
          test_mode)) ;
    mux21 ix1117 (.Y (Result_OUT[23]), .A0 (REG_OUT_23), .A1 (MISR_OUT_23), .S0 (
          test_mode)) ;
    mux21 ix1125 (.Y (Result_OUT[24]), .A0 (REG_OUT_24), .A1 (MISR_OUT_24), .S0 (
          test_mode)) ;
    mux21 ix1133 (.Y (Result_OUT[25]), .A0 (REG_OUT_25), .A1 (MISR_OUT_25), .S0 (
          test_mode)) ;
    mux21 ix1141 (.Y (Result_OUT[26]), .A0 (REG_OUT_26), .A1 (MISR_OUT_26), .S0 (
          test_mode)) ;
    mux21 ix1149 (.Y (Result_OUT[27]), .A0 (REG_OUT_27), .A1 (MISR_OUT_27), .S0 (
          test_mode)) ;
    mux21 ix1157 (.Y (Result_OUT[28]), .A0 (REG_OUT_28), .A1 (MISR_OUT_28), .S0 (
          test_mode)) ;
    mux21 ix1165 (.Y (Result_OUT[29]), .A0 (REG_OUT_29), .A1 (MISR_OUT_29), .S0 (
          test_mode)) ;
    mux21 ix1173 (.Y (Result_OUT[30]), .A0 (REG_OUT_30), .A1 (MISR_OUT_30), .S0 (
          test_mode)) ;
    mux21 ix1181 (.Y (Result_OUT[31]), .A0 (REG_OUT_31), .A1 (MISR_OUT_31), .S0 (
          test_mode)) ;
    inv01 ix1 (.Y (nx0), .A (nx1334)) ;
    inv01 ix1690 (.Y (nx1691), .A (nx1701)) ;
    inv02 ix1692 (.Y (nx1693), .A (nx1705)) ;
    inv02 ix1694 (.Y (nx1695), .A (nx1705)) ;
    inv02 ix1696 (.Y (nx1697), .A (nx1705)) ;
    inv01 ix1698 (.Y (nx1699), .A (nx0)) ;
    inv01 ix1700 (.Y (nx1701), .A (nx0)) ;
    inv02 ix1704 (.Y (nx1705), .A (nx937)) ;
    mux21 ix1312 (.Y (nx1311), .A0 (MISR_EN), .A1 (nx662), .S0 (nx0)) ;
    and04 ix505 (.Y (nx504), .A0 (nx1590), .A1 (nx1331), .A2 (nx1340), .A3 (
          nx1351)) ;
    mux21 ix1292 (.Y (nx1291), .A0 (clk_cnt_30), .A1 (nx484), .S0 (nx1719)) ;
    nor02ii ix459 (.Y (nx981), .A0 (nx1347), .A1 (clk_cnt_28)) ;
    mux21 ix1272 (.Y (nx1271), .A0 (clk_cnt_28), .A1 (nx450), .S0 (nx1719)) ;
    and02 ix1345 (.Y (nx1344), .A0 (nx1340), .A1 (nx1347)) ;
    nor02ii ix427 (.Y (nx979), .A0 (nx1364), .A1 (clk_cnt_26)) ;
    mux21 ix1252 (.Y (nx1251), .A0 (clk_cnt_26), .A1 (nx418), .S0 (nx1719)) ;
    and02 ix1362 (.Y (nx1361), .A0 (nx1357), .A1 (nx1364)) ;
    nor02ii ix395 (.Y (nx975), .A0 (nx1381), .A1 (clk_cnt_24)) ;
    mux21 ix1232 (.Y (nx1231), .A0 (clk_cnt_24), .A1 (nx386), .S0 (nx1719)) ;
    and02 ix1379 (.Y (nx1378), .A0 (nx1374), .A1 (nx1381)) ;
    nor02ii ix363 (.Y (nx972), .A0 (nx1398), .A1 (clk_cnt_22)) ;
    mux21 ix1212 (.Y (nx1211), .A0 (clk_cnt_22), .A1 (nx354), .S0 (nx1719)) ;
    and02 ix1396 (.Y (nx1395), .A0 (nx1391), .A1 (nx1398)) ;
    nor02ii ix331 (.Y (nx969), .A0 (nx1415), .A1 (clk_cnt_20)) ;
    mux21 ix1192 (.Y (nx1191), .A0 (clk_cnt_20), .A1 (nx322), .S0 (nx1719)) ;
    and02 ix1413 (.Y (nx1412), .A0 (nx1408), .A1 (nx1415)) ;
    nor02ii ix299 (.Y (nx965), .A0 (nx1432), .A1 (clk_cnt_18)) ;
    mux21 ix1172 (.Y (nx1171), .A0 (clk_cnt_18), .A1 (nx290), .S0 (nx1719)) ;
    and02 ix1430 (.Y (nx1429), .A0 (nx1425), .A1 (nx1432)) ;
    nor02ii ix267 (.Y (nx963), .A0 (nx1449), .A1 (clk_cnt_16)) ;
    mux21 ix1152 (.Y (nx1151), .A0 (clk_cnt_16), .A1 (nx258), .S0 (nx1719)) ;
    and02 ix1447 (.Y (nx1446), .A0 (nx1442), .A1 (nx1449)) ;
    nor02ii ix235 (.Y (nx959), .A0 (nx1466), .A1 (clk_cnt_14)) ;
    mux21 ix1132 (.Y (nx1131), .A0 (clk_cnt_14), .A1 (nx226), .S0 (nx1719)) ;
    and02 ix1464 (.Y (nx1463), .A0 (nx1459), .A1 (nx1466)) ;
    nor02ii ix203 (.Y (nx956), .A0 (nx1483), .A1 (clk_cnt_12)) ;
    mux21 ix1112 (.Y (nx1111), .A0 (clk_cnt_12), .A1 (nx194), .S0 (nx1719)) ;
    and02 ix1481 (.Y (nx1480), .A0 (nx1476), .A1 (nx1483)) ;
    nor02ii ix171 (.Y (nx953), .A0 (nx1500), .A1 (clk_cnt_10)) ;
    mux21 ix1092 (.Y (nx1091), .A0 (clk_cnt_10), .A1 (nx162), .S0 (nx1721)) ;
    and02 ix1498 (.Y (nx1497), .A0 (nx1493), .A1 (nx1500)) ;
    nor02ii ix139 (.Y (nx949), .A0 (nx1517), .A1 (clk_cnt_8)) ;
    mux21 ix1072 (.Y (nx1071), .A0 (clk_cnt_8), .A1 (nx130), .S0 (nx1721)) ;
    and02 ix1515 (.Y (nx1514), .A0 (nx1510), .A1 (nx1517)) ;
    nor02ii ix107 (.Y (nx947), .A0 (nx1533), .A1 (clk_cnt_6)) ;
    or04 ix1531 (.Y (nx1530), .A0 (nx1711), .A1 (nx1701), .A2 (nx947), .A3 (
         nx1705)) ;
    nor02ii ix93 (.Y (nx1711), .A0 (clk_cnt_6), .A1 (nx1533)) ;
    nor02ii ix75 (.Y (nx943), .A0 (nx1549), .A1 (clk_cnt_4)) ;
    or04 ix1547 (.Y (nx1546), .A0 (nx1713), .A1 (nx1701), .A2 (nx943), .A3 (
         nx1705)) ;
    nor02ii ix61 (.Y (nx1713), .A0 (clk_cnt_4), .A1 (nx1549)) ;
    mux21 ix1002 (.Y (nx1001), .A0 (clk_cnt_1), .A1 (nx18), .S0 (nx1721)) ;
    nor02ii ix19 (.Y (nx18), .A0 (nx1572), .A1 (nx0)) ;
    mux21 ix992 (.Y (nx991), .A0 (clk_cnt_0), .A1 (nx4), .S0 (nx1721)) ;
    nor02ii ix5 (.Y (nx4), .A0 (clk_cnt_0), .A1 (nx0)) ;
    or02 ix1578 (.Y (nx937), .A0 (nx1699), .A1 (nx610)) ;
    and03 ix515 (.Y (nx514), .A0 (nx1374), .A1 (nx1357), .A2 (nx1368)) ;
    and03 ix527 (.Y (nx526), .A0 (nx1402), .A1 (nx1385), .A2 (nx1391)) ;
    and03 ix537 (.Y (nx536), .A0 (nx1425), .A1 (nx1408), .A2 (nx1419)) ;
    and03 ix551 (.Y (nx550), .A0 (nx1453), .A1 (nx1436), .A2 (nx1442)) ;
    and03 ix561 (.Y (nx560), .A0 (nx1476), .A1 (nx1459), .A2 (nx1470)) ;
    and03 ix573 (.Y (nx572), .A0 (nx1504), .A1 (nx1487), .A2 (nx1493)) ;
    ao21 ix583 (.Y (nx582), .A0 (nx1562), .A1 (nx1567), .B0 (nx1553)) ;
    and02 ix589 (.Y (nx588), .A0 (nx1537), .A1 (nx1543)) ;
    and03 ix1300 (.Y (nx1299), .A0 (nx0), .A1 (nx1715), .A2 (nx1721)) ;
    xnor2 ix1612 (.Y (nx1715), .A0 (nx1608), .A1 (nx478)) ;
    nor02ii ix479 (.Y (nx478), .A0 (nx1327), .A1 (clk_cnt_30)) ;
    nor02ii ix1616 (.Y (nx1615), .A0 (nx652), .A1 (nx1608)) ;
    and04 ix653 (.Y (nx652), .A0 (nx1543), .A1 (nx1527), .A2 (nx1537), .A3 (
          nx1717)) ;
    and03 ix1619 (.Y (nx1717), .A0 (nx644), .A1 (nx1553), .A2 (nx610)) ;
    inv01 ix1718 (.Y (nx1719), .A (nx1705)) ;
    inv01 ix1720 (.Y (nx1721), .A (nx1705)) ;
endmodule


module RCFA_32 ( A, B, Cin, Sum, Cout ) ;

    input [31:0]A ;
    input [31:0]B ;
    input Cin ;
    output [31:0]Sum ;
    output Cout ;

    wire nx8, nx10, nx12, nx22, nx28, nx30, nx32, nx42, nx48, nx50, nx52, nx62, 
         nx68, nx70, nx72, nx82, nx88, nx90, nx92, nx102, nx108, nx110, nx112, 
         nx122, nx128, nx130, nx132, nx142, nx148, nx150, nx152, nx162, nx168, 
         nx170, nx172, nx182, nx188, nx190, nx192, nx202, nx208, nx210, nx212, 
         nx222, nx228, nx230, nx232, nx242, nx248, nx250, nx252, nx262, nx268, 
         nx270, nx272, nx282, nx288, nx290, nx292, nx302, nx308, nx310, nx312, 
         nx510, nx514, nx518, nx522, nx526, nx530, nx534, nx538, nx542, nx546, 
         nx550, nx554, nx558, nx562, nx566, nx571, nx573, nx575, nx577, nx580, 
         nx582, nx584, nx586, nx589, nx591, nx593, nx595, nx598, nx600, nx602, 
         nx604, nx607, nx609, nx611, nx613, nx616, nx618, nx620, nx622, nx625, 
         nx627, nx629, nx631, nx634, nx636, nx638, nx640, nx643, nx645, nx647, 
         nx649, nx652, nx654, nx656, nx658, nx661, nx663, nx665, nx667, nx670, 
         nx672, nx674, nx676, nx679, nx681, nx683, nx685, nx688, nx690, nx692, 
         nx694, nx697, nx699, nx701, nx703, nx706;



    ao22 ix321 (.Y (Cout), .A0 (A[31]), .A1 (nx310), .B0 (nx308), .B1 (nx312)) ;
    oai22 ix309 (.Y (nx308), .A0 (nx510), .A1 (nx699), .B0 (nx703), .B1 (nx701)
          ) ;
    aoi22 ix511 (.Y (nx510), .A0 (A[29]), .A1 (nx290), .B0 (nx288), .B1 (nx292)
          ) ;
    oai22 ix289 (.Y (nx288), .A0 (nx514), .A1 (nx690), .B0 (nx694), .B1 (nx692)
          ) ;
    aoi22 ix515 (.Y (nx514), .A0 (A[27]), .A1 (nx270), .B0 (nx268), .B1 (nx272)
          ) ;
    oai22 ix269 (.Y (nx268), .A0 (nx518), .A1 (nx681), .B0 (nx685), .B1 (nx683)
          ) ;
    aoi22 ix519 (.Y (nx518), .A0 (A[25]), .A1 (nx250), .B0 (nx248), .B1 (nx252)
          ) ;
    oai22 ix249 (.Y (nx248), .A0 (nx522), .A1 (nx672), .B0 (nx676), .B1 (nx674)
          ) ;
    aoi22 ix523 (.Y (nx522), .A0 (A[23]), .A1 (nx230), .B0 (nx228), .B1 (nx232)
          ) ;
    oai22 ix229 (.Y (nx228), .A0 (nx526), .A1 (nx663), .B0 (nx667), .B1 (nx665)
          ) ;
    aoi22 ix527 (.Y (nx526), .A0 (A[21]), .A1 (nx210), .B0 (nx208), .B1 (nx212)
          ) ;
    oai22 ix209 (.Y (nx208), .A0 (nx530), .A1 (nx654), .B0 (nx658), .B1 (nx656)
          ) ;
    aoi22 ix531 (.Y (nx530), .A0 (A[19]), .A1 (nx190), .B0 (nx188), .B1 (nx192)
          ) ;
    oai22 ix189 (.Y (nx188), .A0 (nx534), .A1 (nx645), .B0 (nx649), .B1 (nx647)
          ) ;
    aoi22 ix535 (.Y (nx534), .A0 (A[17]), .A1 (nx170), .B0 (nx168), .B1 (nx172)
          ) ;
    oai22 ix169 (.Y (nx168), .A0 (nx538), .A1 (nx636), .B0 (nx640), .B1 (nx638)
          ) ;
    aoi22 ix539 (.Y (nx538), .A0 (A[15]), .A1 (nx150), .B0 (nx148), .B1 (nx152)
          ) ;
    oai22 ix149 (.Y (nx148), .A0 (nx542), .A1 (nx627), .B0 (nx631), .B1 (nx629)
          ) ;
    aoi22 ix543 (.Y (nx542), .A0 (A[13]), .A1 (nx130), .B0 (nx128), .B1 (nx132)
          ) ;
    oai22 ix129 (.Y (nx128), .A0 (nx546), .A1 (nx618), .B0 (nx622), .B1 (nx620)
          ) ;
    aoi22 ix547 (.Y (nx546), .A0 (A[11]), .A1 (nx110), .B0 (nx108), .B1 (nx112)
          ) ;
    oai22 ix109 (.Y (nx108), .A0 (nx550), .A1 (nx609), .B0 (nx613), .B1 (nx611)
          ) ;
    aoi22 ix551 (.Y (nx550), .A0 (A[9]), .A1 (nx90), .B0 (nx88), .B1 (nx92)) ;
    oai22 ix89 (.Y (nx88), .A0 (nx554), .A1 (nx600), .B0 (nx604), .B1 (nx602)) ;
    aoi22 ix555 (.Y (nx554), .A0 (A[7]), .A1 (nx70), .B0 (nx68), .B1 (nx72)) ;
    oai22 ix69 (.Y (nx68), .A0 (nx558), .A1 (nx591), .B0 (nx595), .B1 (nx593)) ;
    aoi22 ix559 (.Y (nx558), .A0 (A[5]), .A1 (nx50), .B0 (nx48), .B1 (nx52)) ;
    oai22 ix49 (.Y (nx48), .A0 (nx562), .A1 (nx582), .B0 (nx586), .B1 (nx584)) ;
    aoi22 ix563 (.Y (nx562), .A0 (A[3]), .A1 (nx30), .B0 (nx28), .B1 (nx32)) ;
    oai22 ix29 (.Y (nx28), .A0 (nx566), .A1 (nx573), .B0 (nx577), .B1 (nx575)) ;
    aoi22 ix567 (.Y (nx566), .A0 (A[1]), .A1 (nx10), .B0 (nx8), .B1 (nx12)) ;
    mux21 ix9 (.Y (nx8), .A0 (Cin), .A1 (A[0]), .S0 (B[0])) ;
    xnor2 ix13 (.Y (nx12), .A0 (A[1]), .A1 (nx571)) ;
    xnor2 ix572 (.Y (nx571), .A0 (B[1]), .A1 (Cin)) ;
    xnor2 ix576 (.Y (nx575), .A0 (B[2]), .A1 (Cin)) ;
    inv01 ix578 (.Y (nx577), .A (A[2])) ;
    xnor2 ix33 (.Y (nx32), .A0 (A[3]), .A1 (nx580)) ;
    xnor2 ix581 (.Y (nx580), .A0 (B[3]), .A1 (Cin)) ;
    xnor2 ix585 (.Y (nx584), .A0 (B[4]), .A1 (Cin)) ;
    inv01 ix587 (.Y (nx586), .A (A[4])) ;
    xnor2 ix53 (.Y (nx52), .A0 (A[5]), .A1 (nx589)) ;
    xnor2 ix590 (.Y (nx589), .A0 (B[5]), .A1 (Cin)) ;
    xnor2 ix594 (.Y (nx593), .A0 (B[6]), .A1 (Cin)) ;
    inv01 ix596 (.Y (nx595), .A (A[6])) ;
    xnor2 ix73 (.Y (nx72), .A0 (A[7]), .A1 (nx598)) ;
    xnor2 ix599 (.Y (nx598), .A0 (B[7]), .A1 (Cin)) ;
    xnor2 ix603 (.Y (nx602), .A0 (B[8]), .A1 (Cin)) ;
    inv01 ix605 (.Y (nx604), .A (A[8])) ;
    xnor2 ix93 (.Y (nx92), .A0 (A[9]), .A1 (nx607)) ;
    xnor2 ix608 (.Y (nx607), .A0 (B[9]), .A1 (Cin)) ;
    xnor2 ix612 (.Y (nx611), .A0 (B[10]), .A1 (Cin)) ;
    inv01 ix614 (.Y (nx613), .A (A[10])) ;
    xnor2 ix113 (.Y (nx112), .A0 (A[11]), .A1 (nx616)) ;
    xnor2 ix617 (.Y (nx616), .A0 (B[11]), .A1 (Cin)) ;
    xnor2 ix621 (.Y (nx620), .A0 (B[12]), .A1 (Cin)) ;
    inv01 ix623 (.Y (nx622), .A (A[12])) ;
    xnor2 ix133 (.Y (nx132), .A0 (A[13]), .A1 (nx625)) ;
    xnor2 ix626 (.Y (nx625), .A0 (B[13]), .A1 (Cin)) ;
    xnor2 ix630 (.Y (nx629), .A0 (B[14]), .A1 (Cin)) ;
    inv01 ix632 (.Y (nx631), .A (A[14])) ;
    xnor2 ix153 (.Y (nx152), .A0 (A[15]), .A1 (nx634)) ;
    xnor2 ix635 (.Y (nx634), .A0 (B[15]), .A1 (Cin)) ;
    xnor2 ix639 (.Y (nx638), .A0 (B[16]), .A1 (Cin)) ;
    inv01 ix641 (.Y (nx640), .A (A[16])) ;
    xnor2 ix173 (.Y (nx172), .A0 (A[17]), .A1 (nx643)) ;
    xnor2 ix644 (.Y (nx643), .A0 (B[17]), .A1 (Cin)) ;
    xnor2 ix648 (.Y (nx647), .A0 (B[18]), .A1 (Cin)) ;
    inv01 ix650 (.Y (nx649), .A (A[18])) ;
    xnor2 ix193 (.Y (nx192), .A0 (A[19]), .A1 (nx652)) ;
    xnor2 ix653 (.Y (nx652), .A0 (B[19]), .A1 (Cin)) ;
    xnor2 ix657 (.Y (nx656), .A0 (B[20]), .A1 (Cin)) ;
    inv01 ix659 (.Y (nx658), .A (A[20])) ;
    xnor2 ix213 (.Y (nx212), .A0 (A[21]), .A1 (nx661)) ;
    xnor2 ix662 (.Y (nx661), .A0 (B[21]), .A1 (Cin)) ;
    xnor2 ix666 (.Y (nx665), .A0 (B[22]), .A1 (Cin)) ;
    inv01 ix668 (.Y (nx667), .A (A[22])) ;
    xnor2 ix233 (.Y (nx232), .A0 (A[23]), .A1 (nx670)) ;
    xnor2 ix671 (.Y (nx670), .A0 (B[23]), .A1 (Cin)) ;
    xnor2 ix675 (.Y (nx674), .A0 (B[24]), .A1 (Cin)) ;
    inv01 ix677 (.Y (nx676), .A (A[24])) ;
    xnor2 ix253 (.Y (nx252), .A0 (A[25]), .A1 (nx679)) ;
    xnor2 ix680 (.Y (nx679), .A0 (B[25]), .A1 (Cin)) ;
    xnor2 ix684 (.Y (nx683), .A0 (B[26]), .A1 (Cin)) ;
    inv01 ix686 (.Y (nx685), .A (A[26])) ;
    xnor2 ix273 (.Y (nx272), .A0 (A[27]), .A1 (nx688)) ;
    xnor2 ix689 (.Y (nx688), .A0 (B[27]), .A1 (Cin)) ;
    xnor2 ix693 (.Y (nx692), .A0 (B[28]), .A1 (Cin)) ;
    inv01 ix695 (.Y (nx694), .A (A[28])) ;
    xnor2 ix293 (.Y (nx292), .A0 (A[29]), .A1 (nx697)) ;
    xnor2 ix698 (.Y (nx697), .A0 (B[29]), .A1 (Cin)) ;
    xnor2 ix702 (.Y (nx701), .A0 (B[30]), .A1 (Cin)) ;
    inv01 ix704 (.Y (nx703), .A (A[30])) ;
    xnor2 ix313 (.Y (nx312), .A0 (A[31]), .A1 (nx706)) ;
    xnor2 ix707 (.Y (nx706), .A0 (B[31]), .A1 (Cin)) ;
    xor2 ix383 (.Y (Sum[0]), .A0 (A[0]), .A1 (B[0])) ;
    xor2 ix381 (.Y (Sum[1]), .A0 (nx8), .A1 (nx12)) ;
    xnor2 ix379 (.Y (Sum[2]), .A0 (nx566), .A1 (nx22)) ;
    xnor2 ix23 (.Y (nx22), .A0 (A[2]), .A1 (nx575)) ;
    xor2 ix377 (.Y (Sum[3]), .A0 (nx28), .A1 (nx32)) ;
    xnor2 ix375 (.Y (Sum[4]), .A0 (nx562), .A1 (nx42)) ;
    xnor2 ix43 (.Y (nx42), .A0 (A[4]), .A1 (nx584)) ;
    xor2 ix373 (.Y (Sum[5]), .A0 (nx48), .A1 (nx52)) ;
    xnor2 ix371 (.Y (Sum[6]), .A0 (nx558), .A1 (nx62)) ;
    xnor2 ix63 (.Y (nx62), .A0 (A[6]), .A1 (nx593)) ;
    xor2 ix369 (.Y (Sum[7]), .A0 (nx68), .A1 (nx72)) ;
    xnor2 ix367 (.Y (Sum[8]), .A0 (nx554), .A1 (nx82)) ;
    xnor2 ix83 (.Y (nx82), .A0 (A[8]), .A1 (nx602)) ;
    xor2 ix365 (.Y (Sum[9]), .A0 (nx88), .A1 (nx92)) ;
    xnor2 ix363 (.Y (Sum[10]), .A0 (nx550), .A1 (nx102)) ;
    xnor2 ix103 (.Y (nx102), .A0 (A[10]), .A1 (nx611)) ;
    xor2 ix361 (.Y (Sum[11]), .A0 (nx108), .A1 (nx112)) ;
    xnor2 ix359 (.Y (Sum[12]), .A0 (nx546), .A1 (nx122)) ;
    xnor2 ix123 (.Y (nx122), .A0 (A[12]), .A1 (nx620)) ;
    xor2 ix357 (.Y (Sum[13]), .A0 (nx128), .A1 (nx132)) ;
    xnor2 ix355 (.Y (Sum[14]), .A0 (nx542), .A1 (nx142)) ;
    xnor2 ix143 (.Y (nx142), .A0 (A[14]), .A1 (nx629)) ;
    xor2 ix353 (.Y (Sum[15]), .A0 (nx148), .A1 (nx152)) ;
    xnor2 ix351 (.Y (Sum[16]), .A0 (nx538), .A1 (nx162)) ;
    xnor2 ix163 (.Y (nx162), .A0 (A[16]), .A1 (nx638)) ;
    xor2 ix349 (.Y (Sum[17]), .A0 (nx168), .A1 (nx172)) ;
    xnor2 ix347 (.Y (Sum[18]), .A0 (nx534), .A1 (nx182)) ;
    xnor2 ix183 (.Y (nx182), .A0 (A[18]), .A1 (nx647)) ;
    xor2 ix345 (.Y (Sum[19]), .A0 (nx188), .A1 (nx192)) ;
    xnor2 ix343 (.Y (Sum[20]), .A0 (nx530), .A1 (nx202)) ;
    xnor2 ix203 (.Y (nx202), .A0 (A[20]), .A1 (nx656)) ;
    xor2 ix341 (.Y (Sum[21]), .A0 (nx208), .A1 (nx212)) ;
    xnor2 ix339 (.Y (Sum[22]), .A0 (nx526), .A1 (nx222)) ;
    xnor2 ix223 (.Y (nx222), .A0 (A[22]), .A1 (nx665)) ;
    xor2 ix337 (.Y (Sum[23]), .A0 (nx228), .A1 (nx232)) ;
    xnor2 ix335 (.Y (Sum[24]), .A0 (nx522), .A1 (nx242)) ;
    xnor2 ix243 (.Y (nx242), .A0 (A[24]), .A1 (nx674)) ;
    xor2 ix333 (.Y (Sum[25]), .A0 (nx248), .A1 (nx252)) ;
    xnor2 ix331 (.Y (Sum[26]), .A0 (nx518), .A1 (nx262)) ;
    xnor2 ix263 (.Y (nx262), .A0 (A[26]), .A1 (nx683)) ;
    xor2 ix329 (.Y (Sum[27]), .A0 (nx268), .A1 (nx272)) ;
    xnor2 ix327 (.Y (Sum[28]), .A0 (nx514), .A1 (nx282)) ;
    xnor2 ix283 (.Y (nx282), .A0 (A[28]), .A1 (nx692)) ;
    xor2 ix325 (.Y (Sum[29]), .A0 (nx288), .A1 (nx292)) ;
    xnor2 ix323 (.Y (Sum[30]), .A0 (nx510), .A1 (nx302)) ;
    xnor2 ix303 (.Y (nx302), .A0 (A[30]), .A1 (nx701)) ;
    xor2 ix315 (.Y (Sum[31]), .A0 (nx308), .A1 (nx312)) ;
    inv01 ix311 (.Y (nx310), .A (nx706)) ;
    inv01 ix700 (.Y (nx699), .A (nx302)) ;
    inv01 ix291 (.Y (nx290), .A (nx697)) ;
    inv01 ix691 (.Y (nx690), .A (nx282)) ;
    inv01 ix271 (.Y (nx270), .A (nx688)) ;
    inv01 ix682 (.Y (nx681), .A (nx262)) ;
    inv01 ix251 (.Y (nx250), .A (nx679)) ;
    inv01 ix673 (.Y (nx672), .A (nx242)) ;
    inv01 ix231 (.Y (nx230), .A (nx670)) ;
    inv01 ix664 (.Y (nx663), .A (nx222)) ;
    inv01 ix211 (.Y (nx210), .A (nx661)) ;
    inv01 ix655 (.Y (nx654), .A (nx202)) ;
    inv01 ix191 (.Y (nx190), .A (nx652)) ;
    inv01 ix646 (.Y (nx645), .A (nx182)) ;
    inv01 ix171 (.Y (nx170), .A (nx643)) ;
    inv01 ix637 (.Y (nx636), .A (nx162)) ;
    inv01 ix151 (.Y (nx150), .A (nx634)) ;
    inv01 ix628 (.Y (nx627), .A (nx142)) ;
    inv01 ix131 (.Y (nx130), .A (nx625)) ;
    inv01 ix619 (.Y (nx618), .A (nx122)) ;
    inv01 ix111 (.Y (nx110), .A (nx616)) ;
    inv01 ix610 (.Y (nx609), .A (nx102)) ;
    inv01 ix91 (.Y (nx90), .A (nx607)) ;
    inv01 ix601 (.Y (nx600), .A (nx82)) ;
    inv01 ix71 (.Y (nx70), .A (nx598)) ;
    inv01 ix592 (.Y (nx591), .A (nx62)) ;
    inv01 ix51 (.Y (nx50), .A (nx589)) ;
    inv01 ix583 (.Y (nx582), .A (nx42)) ;
    inv01 ix31 (.Y (nx30), .A (nx580)) ;
    inv01 ix574 (.Y (nx573), .A (nx22)) ;
    inv01 ix11 (.Y (nx10), .A (nx571)) ;
endmodule


module MISR ( clk, rst, enable, mult_result, signature ) ;

    input clk ;
    input rst ;
    input enable ;
    input [31:0]mult_result ;
    output [31:0]signature ;

    wire zeroth_in, nx12, nx22, nx34, nx44, nx54, nx64, nx76, nx88, nx98, nx108, 
         nx118, nx128, nx138, nx148, nx158, nx168, nx178, nx188, nx198, nx208, 
         nx218, nx228, nx238, nx248, nx258, nx268, nx278, nx288, nx298, nx308, 
         nx318, nx328, nx836, nx846, nx856, nx866, nx876, nx886, nx896, nx906, 
         nx916, nx926, nx936, nx946, nx956, nx966, nx976, nx986, nx996, nx1006, 
         nx1016, nx1026, nx1036, nx1046, nx1056, nx1066, nx1076, nx1086, nx1096, 
         nx1106, nx1116, nx1126, nx1136, nx1146, nx1156, nx1168, nx1170, nx1245, 
         nx1250, nx1264, nx1272, nx1276, nx1315, nx1317, nx1323, nx1325, nx1327, 
         nx1329;
    wire [31:0] \$dummy ;




    dff reg_MISR_REG_0 (.Q (signature[0]), .QB (\$dummy [0]), .D (nx1156), .CLK (
        clk)) ;
    ao221 ix1157 (.Y (nx1156), .A0 (signature[0]), .A1 (nx1315), .B0 (nx328), .B1 (
          nx1329), .C0 (nx1170)) ;
    inv01 ix1171 (.Y (nx1170), .A (rst)) ;
    xor2 ix329 (.Y (nx328), .A0 (mult_result[0]), .A1 (signature[1])) ;
    dff reg_MISR_REG_1 (.Q (signature[1]), .QB (\$dummy [1]), .D (nx1146), .CLK (
        clk)) ;
    ao32 ix1147 (.Y (nx1146), .A0 (rst), .A1 (nx318), .A2 (nx1329), .B0 (
         signature[1]), .B1 (nx1168)) ;
    xor2 ix319 (.Y (nx318), .A0 (mult_result[1]), .A1 (signature[2])) ;
    dff reg_MISR_REG_2 (.Q (signature[2]), .QB (\$dummy [2]), .D (nx1136), .CLK (
        clk)) ;
    ao32 ix1137 (.Y (nx1136), .A0 (rst), .A1 (nx308), .A2 (nx1329), .B0 (
         signature[2]), .B1 (nx1168)) ;
    xor2 ix309 (.Y (nx308), .A0 (mult_result[2]), .A1 (signature[3])) ;
    dff reg_MISR_REG_3 (.Q (signature[3]), .QB (\$dummy [3]), .D (nx1126), .CLK (
        clk)) ;
    ao32 ix1127 (.Y (nx1126), .A0 (rst), .A1 (nx298), .A2 (nx1327), .B0 (
         signature[3]), .B1 (nx1168)) ;
    xor2 ix299 (.Y (nx298), .A0 (mult_result[3]), .A1 (signature[4])) ;
    dff reg_MISR_REG_4 (.Q (signature[4]), .QB (\$dummy [4]), .D (nx1116), .CLK (
        clk)) ;
    ao32 ix1117 (.Y (nx1116), .A0 (rst), .A1 (nx288), .A2 (nx1327), .B0 (
         signature[4]), .B1 (nx1317)) ;
    xor2 ix289 (.Y (nx288), .A0 (mult_result[4]), .A1 (signature[5])) ;
    dff reg_MISR_REG_5 (.Q (signature[5]), .QB (\$dummy [5]), .D (nx1106), .CLK (
        clk)) ;
    ao32 ix1107 (.Y (nx1106), .A0 (rst), .A1 (nx278), .A2 (nx1327), .B0 (
         signature[5]), .B1 (nx1317)) ;
    xor2 ix279 (.Y (nx278), .A0 (mult_result[5]), .A1 (signature[6])) ;
    dff reg_MISR_REG_6 (.Q (signature[6]), .QB (\$dummy [6]), .D (nx1096), .CLK (
        clk)) ;
    ao32 ix1097 (.Y (nx1096), .A0 (rst), .A1 (nx268), .A2 (nx1327), .B0 (
         signature[6]), .B1 (nx1317)) ;
    xor2 ix269 (.Y (nx268), .A0 (mult_result[6]), .A1 (signature[7])) ;
    dff reg_MISR_REG_7 (.Q (signature[7]), .QB (\$dummy [7]), .D (nx1086), .CLK (
        clk)) ;
    ao32 ix1087 (.Y (nx1086), .A0 (rst), .A1 (nx258), .A2 (nx1327), .B0 (
         signature[7]), .B1 (nx1317)) ;
    xor2 ix259 (.Y (nx258), .A0 (mult_result[7]), .A1 (signature[8])) ;
    dff reg_MISR_REG_8 (.Q (signature[8]), .QB (\$dummy [8]), .D (nx1076), .CLK (
        clk)) ;
    ao32 ix1077 (.Y (nx1076), .A0 (rst), .A1 (nx248), .A2 (nx1327), .B0 (
         signature[8]), .B1 (nx1317)) ;
    xor2 ix249 (.Y (nx248), .A0 (mult_result[8]), .A1 (signature[9])) ;
    dff reg_MISR_REG_9 (.Q (signature[9]), .QB (\$dummy [9]), .D (nx1066), .CLK (
        clk)) ;
    ao32 ix1067 (.Y (nx1066), .A0 (rst), .A1 (nx238), .A2 (nx1327), .B0 (
         signature[9]), .B1 (nx1317)) ;
    xor2 ix239 (.Y (nx238), .A0 (mult_result[9]), .A1 (signature[10])) ;
    dff reg_MISR_REG_10 (.Q (signature[10]), .QB (\$dummy [10]), .D (nx1056), .CLK (
        clk)) ;
    ao32 ix1057 (.Y (nx1056), .A0 (rst), .A1 (nx228), .A2 (nx1327), .B0 (
         signature[10]), .B1 (nx1317)) ;
    xor2 ix229 (.Y (nx228), .A0 (mult_result[10]), .A1 (signature[11])) ;
    dff reg_MISR_REG_11 (.Q (signature[11]), .QB (\$dummy [11]), .D (nx1046), .CLK (
        clk)) ;
    ao32 ix1047 (.Y (nx1046), .A0 (rst), .A1 (nx218), .A2 (nx1327), .B0 (
         signature[11]), .B1 (nx1317)) ;
    xor2 ix219 (.Y (nx218), .A0 (mult_result[11]), .A1 (signature[12])) ;
    dff reg_MISR_REG_12 (.Q (signature[12]), .QB (\$dummy [12]), .D (nx1036), .CLK (
        clk)) ;
    ao32 ix1037 (.Y (nx1036), .A0 (rst), .A1 (nx208), .A2 (nx1327), .B0 (
         signature[12]), .B1 (nx1317)) ;
    xor2 ix209 (.Y (nx208), .A0 (mult_result[12]), .A1 (signature[13])) ;
    dff reg_MISR_REG_13 (.Q (signature[13]), .QB (\$dummy [13]), .D (nx1026), .CLK (
        clk)) ;
    ao32 ix1027 (.Y (nx1026), .A0 (rst), .A1 (nx198), .A2 (nx1327), .B0 (
         signature[13]), .B1 (nx1317)) ;
    xor2 ix199 (.Y (nx198), .A0 (mult_result[13]), .A1 (signature[14])) ;
    dff reg_MISR_REG_14 (.Q (signature[14]), .QB (\$dummy [14]), .D (nx1016), .CLK (
        clk)) ;
    ao32 ix1017 (.Y (nx1016), .A0 (rst), .A1 (nx188), .A2 (nx1327), .B0 (
         signature[14]), .B1 (nx1317)) ;
    xor2 ix189 (.Y (nx188), .A0 (mult_result[14]), .A1 (signature[15])) ;
    dff reg_MISR_REG_15 (.Q (signature[15]), .QB (\$dummy [15]), .D (nx1006), .CLK (
        clk)) ;
    ao32 ix1007 (.Y (nx1006), .A0 (rst), .A1 (nx178), .A2 (nx1327), .B0 (
         signature[15]), .B1 (nx1317)) ;
    xor2 ix179 (.Y (nx178), .A0 (mult_result[15]), .A1 (signature[16])) ;
    dff reg_MISR_REG_16 (.Q (signature[16]), .QB (\$dummy [16]), .D (nx996), .CLK (
        clk)) ;
    ao32 ix997 (.Y (nx996), .A0 (rst), .A1 (nx168), .A2 (nx1327), .B0 (
         signature[16]), .B1 (nx1317)) ;
    xor2 ix169 (.Y (nx168), .A0 (mult_result[16]), .A1 (signature[17])) ;
    dff reg_MISR_REG_17 (.Q (signature[17]), .QB (\$dummy [17]), .D (nx986), .CLK (
        clk)) ;
    ao32 ix987 (.Y (nx986), .A0 (rst), .A1 (nx158), .A2 (nx1327), .B0 (
         signature[17]), .B1 (nx1317)) ;
    xor2 ix159 (.Y (nx158), .A0 (mult_result[17]), .A1 (signature[18])) ;
    dff reg_MISR_REG_18 (.Q (signature[18]), .QB (\$dummy [18]), .D (nx976), .CLK (
        clk)) ;
    ao32 ix977 (.Y (nx976), .A0 (rst), .A1 (nx148), .A2 (nx1325), .B0 (
         signature[18]), .B1 (nx1317)) ;
    xor2 ix149 (.Y (nx148), .A0 (mult_result[18]), .A1 (signature[19])) ;
    dff reg_MISR_REG_19 (.Q (signature[19]), .QB (\$dummy [19]), .D (nx966), .CLK (
        clk)) ;
    ao32 ix967 (.Y (nx966), .A0 (rst), .A1 (nx138), .A2 (nx1325), .B0 (
         signature[19]), .B1 (nx1315)) ;
    xor2 ix139 (.Y (nx138), .A0 (mult_result[19]), .A1 (signature[20])) ;
    dff reg_MISR_REG_20 (.Q (signature[20]), .QB (\$dummy [20]), .D (nx956), .CLK (
        clk)) ;
    ao32 ix957 (.Y (nx956), .A0 (rst), .A1 (nx128), .A2 (nx1325), .B0 (
         signature[20]), .B1 (nx1315)) ;
    xor2 ix129 (.Y (nx128), .A0 (mult_result[20]), .A1 (signature[21])) ;
    dff reg_MISR_REG_21 (.Q (signature[21]), .QB (\$dummy [21]), .D (nx946), .CLK (
        clk)) ;
    ao32 ix947 (.Y (nx946), .A0 (rst), .A1 (nx118), .A2 (nx1325), .B0 (
         signature[21]), .B1 (nx1315)) ;
    xor2 ix119 (.Y (nx118), .A0 (mult_result[21]), .A1 (signature[22])) ;
    dff reg_MISR_REG_22 (.Q (signature[22]), .QB (\$dummy [22]), .D (nx936), .CLK (
        clk)) ;
    ao32 ix937 (.Y (nx936), .A0 (rst), .A1 (nx108), .A2 (nx1325), .B0 (
         signature[22]), .B1 (nx1315)) ;
    xor2 ix109 (.Y (nx108), .A0 (mult_result[22]), .A1 (signature[23])) ;
    dff reg_MISR_REG_23 (.Q (signature[23]), .QB (\$dummy [23]), .D (nx926), .CLK (
        clk)) ;
    ao32 ix927 (.Y (nx926), .A0 (rst), .A1 (nx98), .A2 (nx1325), .B0 (
         signature[23]), .B1 (nx1315)) ;
    xor2 ix99 (.Y (nx98), .A0 (mult_result[23]), .A1 (signature[24])) ;
    dff reg_MISR_REG_24 (.Q (signature[24]), .QB (\$dummy [24]), .D (nx916), .CLK (
        clk)) ;
    ao32 ix917 (.Y (nx916), .A0 (rst), .A1 (nx88), .A2 (nx1325), .B0 (
         signature[24]), .B1 (nx1315)) ;
    xnor2 ix1246 (.Y (nx1245), .A0 (mult_result[24]), .A1 (signature[25])) ;
    dff reg_MISR_REG_25 (.Q (signature[25]), .QB (\$dummy [25]), .D (nx906), .CLK (
        clk)) ;
    ao32 ix907 (.Y (nx906), .A0 (rst), .A1 (nx76), .A2 (nx1325), .B0 (
         signature[25]), .B1 (nx1315)) ;
    xnor2 ix1251 (.Y (nx1250), .A0 (mult_result[25]), .A1 (signature[26])) ;
    dff reg_MISR_REG_26 (.Q (signature[26]), .QB (\$dummy [26]), .D (nx896), .CLK (
        clk)) ;
    ao32 ix897 (.Y (nx896), .A0 (rst), .A1 (nx64), .A2 (nx1325), .B0 (
         signature[26]), .B1 (nx1315)) ;
    xor2 ix65 (.Y (nx64), .A0 (mult_result[26]), .A1 (signature[27])) ;
    dff reg_MISR_REG_27 (.Q (signature[27]), .QB (\$dummy [27]), .D (nx886), .CLK (
        clk)) ;
    ao32 ix887 (.Y (nx886), .A0 (rst), .A1 (nx54), .A2 (nx1325), .B0 (
         signature[27]), .B1 (nx1315)) ;
    xor2 ix55 (.Y (nx54), .A0 (mult_result[27]), .A1 (signature[28])) ;
    dff reg_MISR_REG_28 (.Q (signature[28]), .QB (\$dummy [28]), .D (nx876), .CLK (
        clk)) ;
    ao32 ix877 (.Y (nx876), .A0 (rst), .A1 (nx44), .A2 (nx1325), .B0 (
         signature[28]), .B1 (nx1315)) ;
    xor2 ix45 (.Y (nx44), .A0 (mult_result[28]), .A1 (signature[29])) ;
    dff reg_MISR_REG_29 (.Q (signature[29]), .QB (\$dummy [29]), .D (nx866), .CLK (
        clk)) ;
    ao32 ix867 (.Y (nx866), .A0 (rst), .A1 (nx34), .A2 (nx1325), .B0 (
         signature[29]), .B1 (nx1315)) ;
    xnor2 ix1265 (.Y (nx1264), .A0 (mult_result[29]), .A1 (signature[30])) ;
    dff reg_MISR_REG_30 (.Q (signature[30]), .QB (\$dummy [30]), .D (nx856), .CLK (
        clk)) ;
    ao32 ix857 (.Y (nx856), .A0 (rst), .A1 (nx22), .A2 (nx1325), .B0 (
         signature[30]), .B1 (nx1315)) ;
    xor2 ix23 (.Y (nx22), .A0 (mult_result[30]), .A1 (signature[31])) ;
    dff reg_MISR_REG_31 (.Q (signature[31]), .QB (\$dummy [31]), .D (nx846), .CLK (
        clk)) ;
    ao32 ix847 (.Y (nx846), .A0 (rst), .A1 (nx12), .A2 (nx1325), .B0 (
         signature[31]), .B1 (nx1315)) ;
    mux21 ix837 (.Y (nx836), .A0 (signature[0]), .A1 (zeroth_in), .S0 (nx1276)
          ) ;
    dff reg_zeroth_in (.Q (zeroth_in), .QB (nx1272), .D (nx836), .CLK (clk)) ;
    nand02 ix1277 (.Y (nx1276), .A0 (nx1325), .A1 (rst)) ;
    nor02ii ix1169 (.Y (nx1168), .A0 (nx1329), .A1 (rst)) ;
    xor2 ix89 (.Y (nx88), .A0 (nx1245), .A1 (nx1272)) ;
    xor2 ix77 (.Y (nx76), .A0 (nx1250), .A1 (nx1272)) ;
    xor2 ix35 (.Y (nx34), .A0 (nx1264), .A1 (nx1272)) ;
    xor2 ix13 (.Y (nx12), .A0 (mult_result[31]), .A1 (zeroth_in)) ;
    nor02ii ix1314 (.Y (nx1315), .A0 (nx1329), .A1 (rst)) ;
    nor02ii ix1316 (.Y (nx1317), .A0 (nx1329), .A1 (rst)) ;
    inv01 ix1322 (.Y (nx1323), .A (enable)) ;
    inv01 ix1324 (.Y (nx1325), .A (nx1323)) ;
    inv01 ix1326 (.Y (nx1327), .A (nx1323)) ;
    inv01 ix1328 (.Y (nx1329), .A (nx1323)) ;
endmodule


module LFSR ( clk, rst, enable, bit_pattern ) ;

    input clk ;
    input rst ;
    input enable ;
    output [31:0]bit_pattern ;

    wire zeroth_in, nx38, nx72, nx82, nx740, nx750, nx760, nx770, nx780, nx790, 
         nx800, nx810, nx820, nx830, nx840, nx850, nx860, nx870, nx880, nx890, 
         nx900, nx910, nx920, nx930, nx940, nx950, nx960, nx970, nx980, nx990, 
         nx1000, nx1010, nx1020, nx1030, nx1040, nx1050, nx1060, nx1139, nx1144, 
         nx1183, nx1185, nx1187, nx1189;
    wire [32:0] \$dummy ;




    dff reg_LFSR_REG_0 (.Q (bit_pattern[0]), .QB (\$dummy [0]), .D (nx740), .CLK (
        clk)) ;
    ao221 ix741 (.Y (nx740), .A0 (bit_pattern[1]), .A1 (enable), .B0 (
          bit_pattern[0]), .B1 (nx1189), .C0 (nx1144)) ;
    dff reg_LFSR_REG_1 (.Q (bit_pattern[1]), .QB (\$dummy [1]), .D (nx1060), .CLK (
        clk)) ;
    ao32 ix1061 (.Y (nx1060), .A0 (rst), .A1 (bit_pattern[2]), .A2 (enable), .B0 (
         bit_pattern[1]), .B1 (nx1189)) ;
    dff reg_LFSR_REG_2 (.Q (bit_pattern[2]), .QB (\$dummy [2]), .D (nx1050), .CLK (
        clk)) ;
    ao32 ix1051 (.Y (nx1050), .A0 (rst), .A1 (bit_pattern[3]), .A2 (enable), .B0 (
         bit_pattern[2]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_3 (.Q (bit_pattern[3]), .QB (\$dummy [3]), .D (nx1040), .CLK (
        clk)) ;
    ao32 ix1041 (.Y (nx1040), .A0 (rst), .A1 (bit_pattern[4]), .A2 (enable), .B0 (
         bit_pattern[3]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_4 (.Q (bit_pattern[4]), .QB (\$dummy [4]), .D (nx1030), .CLK (
        clk)) ;
    ao32 ix1031 (.Y (nx1030), .A0 (rst), .A1 (bit_pattern[5]), .A2 (enable), .B0 (
         bit_pattern[4]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_5 (.Q (bit_pattern[5]), .QB (\$dummy [5]), .D (nx1020), .CLK (
        clk)) ;
    ao32 ix1021 (.Y (nx1020), .A0 (rst), .A1 (bit_pattern[6]), .A2 (enable), .B0 (
         bit_pattern[5]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_6 (.Q (bit_pattern[6]), .QB (\$dummy [6]), .D (nx1010), .CLK (
        clk)) ;
    ao32 ix1011 (.Y (nx1010), .A0 (rst), .A1 (bit_pattern[7]), .A2 (enable), .B0 (
         bit_pattern[6]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_7 (.Q (bit_pattern[7]), .QB (\$dummy [7]), .D (nx1000), .CLK (
        clk)) ;
    ao32 ix1001 (.Y (nx1000), .A0 (rst), .A1 (bit_pattern[8]), .A2 (enable), .B0 (
         bit_pattern[7]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_8 (.Q (bit_pattern[8]), .QB (\$dummy [8]), .D (nx990), .CLK (
        clk)) ;
    ao32 ix991 (.Y (nx990), .A0 (rst), .A1 (bit_pattern[9]), .A2 (enable), .B0 (
         bit_pattern[8]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_9 (.Q (bit_pattern[9]), .QB (\$dummy [9]), .D (nx980), .CLK (
        clk)) ;
    ao32 ix981 (.Y (nx980), .A0 (rst), .A1 (bit_pattern[10]), .A2 (enable), .B0 (
         bit_pattern[9]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_10 (.Q (bit_pattern[10]), .QB (\$dummy [10]), .D (nx970), .CLK (
        clk)) ;
    ao32 ix971 (.Y (nx970), .A0 (rst), .A1 (bit_pattern[11]), .A2 (enable), .B0 (
         bit_pattern[10]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_11 (.Q (bit_pattern[11]), .QB (\$dummy [11]), .D (nx960), .CLK (
        clk)) ;
    ao32 ix961 (.Y (nx960), .A0 (rst), .A1 (bit_pattern[12]), .A2 (enable), .B0 (
         bit_pattern[11]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_12 (.Q (bit_pattern[12]), .QB (\$dummy [12]), .D (nx950), .CLK (
        clk)) ;
    ao32 ix951 (.Y (nx950), .A0 (rst), .A1 (bit_pattern[13]), .A2 (enable), .B0 (
         bit_pattern[12]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_13 (.Q (bit_pattern[13]), .QB (\$dummy [13]), .D (nx940), .CLK (
        clk)) ;
    ao32 ix941 (.Y (nx940), .A0 (rst), .A1 (bit_pattern[14]), .A2 (enable), .B0 (
         bit_pattern[13]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_14 (.Q (bit_pattern[14]), .QB (\$dummy [14]), .D (nx930), .CLK (
        clk)) ;
    ao32 ix931 (.Y (nx930), .A0 (rst), .A1 (bit_pattern[15]), .A2 (enable), .B0 (
         bit_pattern[14]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_15 (.Q (bit_pattern[15]), .QB (\$dummy [15]), .D (nx920), .CLK (
        clk)) ;
    ao32 ix921 (.Y (nx920), .A0 (rst), .A1 (bit_pattern[16]), .A2 (enable), .B0 (
         bit_pattern[15]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_16 (.Q (bit_pattern[16]), .QB (\$dummy [16]), .D (nx910), .CLK (
        clk)) ;
    ao32 ix911 (.Y (nx910), .A0 (rst), .A1 (bit_pattern[17]), .A2 (enable), .B0 (
         bit_pattern[16]), .B1 (nx1187)) ;
    dff reg_LFSR_REG_17 (.Q (bit_pattern[17]), .QB (\$dummy [17]), .D (nx900), .CLK (
        clk)) ;
    ao32 ix901 (.Y (nx900), .A0 (rst), .A1 (bit_pattern[18]), .A2 (enable), .B0 (
         bit_pattern[17]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_18 (.Q (bit_pattern[18]), .QB (\$dummy [18]), .D (nx890), .CLK (
        clk)) ;
    ao32 ix891 (.Y (nx890), .A0 (rst), .A1 (bit_pattern[19]), .A2 (enable), .B0 (
         bit_pattern[18]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_19 (.Q (bit_pattern[19]), .QB (\$dummy [19]), .D (nx880), .CLK (
        clk)) ;
    ao32 ix881 (.Y (nx880), .A0 (rst), .A1 (bit_pattern[20]), .A2 (enable), .B0 (
         bit_pattern[19]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_20 (.Q (bit_pattern[20]), .QB (\$dummy [20]), .D (nx870), .CLK (
        clk)) ;
    ao32 ix871 (.Y (nx870), .A0 (rst), .A1 (bit_pattern[21]), .A2 (enable), .B0 (
         bit_pattern[20]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_21 (.Q (bit_pattern[21]), .QB (\$dummy [21]), .D (nx860), .CLK (
        clk)) ;
    ao32 ix861 (.Y (nx860), .A0 (rst), .A1 (bit_pattern[22]), .A2 (enable), .B0 (
         bit_pattern[21]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_22 (.Q (bit_pattern[22]), .QB (\$dummy [22]), .D (nx850), .CLK (
        clk)) ;
    ao32 ix851 (.Y (nx850), .A0 (rst), .A1 (bit_pattern[23]), .A2 (enable), .B0 (
         bit_pattern[22]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_23 (.Q (bit_pattern[23]), .QB (\$dummy [23]), .D (nx840), .CLK (
        clk)) ;
    ao32 ix841 (.Y (nx840), .A0 (rst), .A1 (bit_pattern[24]), .A2 (enable), .B0 (
         bit_pattern[23]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_24 (.Q (bit_pattern[24]), .QB (\$dummy [24]), .D (nx830), .CLK (
        clk)) ;
    ao32 ix831 (.Y (nx830), .A0 (rst), .A1 (nx82), .A2 (enable), .B0 (
         bit_pattern[24]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_25 (.Q (bit_pattern[25]), .QB (\$dummy [25]), .D (nx820), .CLK (
        clk)) ;
    ao32 ix821 (.Y (nx820), .A0 (rst), .A1 (nx72), .A2 (enable), .B0 (
         bit_pattern[25]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_26 (.Q (bit_pattern[26]), .QB (\$dummy [26]), .D (nx810), .CLK (
        clk)) ;
    ao32 ix811 (.Y (nx810), .A0 (rst), .A1 (bit_pattern[27]), .A2 (enable), .B0 (
         bit_pattern[26]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_27 (.Q (bit_pattern[27]), .QB (\$dummy [27]), .D (nx800), .CLK (
        clk)) ;
    ao32 ix801 (.Y (nx800), .A0 (rst), .A1 (bit_pattern[28]), .A2 (enable), .B0 (
         bit_pattern[27]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_28 (.Q (bit_pattern[28]), .QB (\$dummy [28]), .D (nx790), .CLK (
        clk)) ;
    ao32 ix791 (.Y (nx790), .A0 (rst), .A1 (bit_pattern[29]), .A2 (enable), .B0 (
         bit_pattern[28]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_29 (.Q (bit_pattern[29]), .QB (\$dummy [29]), .D (nx780), .CLK (
        clk)) ;
    ao32 ix781 (.Y (nx780), .A0 (rst), .A1 (nx38), .A2 (enable), .B0 (
         bit_pattern[29]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_30 (.Q (bit_pattern[30]), .QB (\$dummy [30]), .D (nx770), .CLK (
        clk)) ;
    ao32 ix771 (.Y (nx770), .A0 (rst), .A1 (bit_pattern[31]), .A2 (enable), .B0 (
         bit_pattern[30]), .B1 (nx1185)) ;
    dff reg_LFSR_REG_31 (.Q (bit_pattern[31]), .QB (\$dummy [31]), .D (nx760), .CLK (
        clk)) ;
    ao32 ix761 (.Y (nx760), .A0 (rst), .A1 (zeroth_in), .A2 (enable), .B0 (
         bit_pattern[31]), .B1 (nx1185)) ;
    dff reg_zeroth_in (.Q (zeroth_in), .QB (\$dummy [32]), .D (nx750), .CLK (clk
        )) ;
    mux21 ix751 (.Y (nx750), .A0 (bit_pattern[0]), .A1 (zeroth_in), .S0 (nx1139)
          ) ;
    nand02 ix1140 (.Y (nx1139), .A0 (enable), .A1 (rst)) ;
    inv01 ix1145 (.Y (nx1144), .A (rst)) ;
    inv01 ix1184 (.Y (nx1185), .A (nx1183)) ;
    inv01 ix1186 (.Y (nx1187), .A (nx1183)) ;
    inv01 ix1188 (.Y (nx1189), .A (nx1183)) ;
    xor2 ix83 (.Y (nx82), .A0 (bit_pattern[25]), .A1 (zeroth_in)) ;
    xor2 ix73 (.Y (nx72), .A0 (bit_pattern[26]), .A1 (zeroth_in)) ;
    xor2 ix39 (.Y (nx38), .A0 (bit_pattern[30]), .A1 (zeroth_in)) ;
    or02 ix1143 (.Y (nx1183), .A0 (nx1144), .A1 (enable)) ;
endmodule


module RegisterN_32 ( clk, reset, enable, \input , \output  ) ;

    input clk ;
    input reset ;
    input enable ;
    input [31:0]\input  ;
    output [31:0]\output  ;

    wire NOT_reset, nx422, nx432, nx442, nx452, nx462, nx472, nx482, nx492, 
         nx502, nx512, nx522, nx532, nx542, nx552, nx562, nx572, nx582, nx592, 
         nx602, nx612, nx622, nx632, nx642, nx652, nx662, nx672, nx682, nx692, 
         nx702, nx712, nx722, nx732, nx845, nx847;
    wire [31:0] \$dummy ;




    dffr reg_output_0 (.Q (\output [0]), .QB (\$dummy [0]), .D (nx422), .CLK (
         clk), .R (nx845)) ;
    mux21 ix423 (.Y (nx422), .A0 (\output [0]), .A1 (\input [0]), .S0 (enable)
          ) ;
    inv01 ix745 (.Y (NOT_reset), .A (reset)) ;
    dffr reg_output_1 (.Q (\output [1]), .QB (\$dummy [1]), .D (nx432), .CLK (
         clk), .R (nx845)) ;
    mux21 ix433 (.Y (nx432), .A0 (\output [1]), .A1 (\input [1]), .S0 (enable)
          ) ;
    dffr reg_output_2 (.Q (\output [2]), .QB (\$dummy [2]), .D (nx442), .CLK (
         clk), .R (nx845)) ;
    mux21 ix443 (.Y (nx442), .A0 (\output [2]), .A1 (\input [2]), .S0 (enable)
          ) ;
    dffr reg_output_3 (.Q (\output [3]), .QB (\$dummy [3]), .D (nx452), .CLK (
         clk), .R (nx845)) ;
    mux21 ix453 (.Y (nx452), .A0 (\output [3]), .A1 (\input [3]), .S0 (enable)
          ) ;
    dffr reg_output_4 (.Q (\output [4]), .QB (\$dummy [4]), .D (nx462), .CLK (
         clk), .R (nx845)) ;
    mux21 ix463 (.Y (nx462), .A0 (\output [4]), .A1 (\input [4]), .S0 (enable)
          ) ;
    dffr reg_output_5 (.Q (\output [5]), .QB (\$dummy [5]), .D (nx472), .CLK (
         clk), .R (nx845)) ;
    mux21 ix473 (.Y (nx472), .A0 (\output [5]), .A1 (\input [5]), .S0 (enable)
          ) ;
    dffr reg_output_6 (.Q (\output [6]), .QB (\$dummy [6]), .D (nx482), .CLK (
         clk), .R (nx845)) ;
    mux21 ix483 (.Y (nx482), .A0 (\output [6]), .A1 (\input [6]), .S0 (enable)
          ) ;
    dffr reg_output_7 (.Q (\output [7]), .QB (\$dummy [7]), .D (nx492), .CLK (
         clk), .R (nx845)) ;
    mux21 ix493 (.Y (nx492), .A0 (\output [7]), .A1 (\input [7]), .S0 (enable)
          ) ;
    dffr reg_output_8 (.Q (\output [8]), .QB (\$dummy [8]), .D (nx502), .CLK (
         clk), .R (nx845)) ;
    mux21 ix503 (.Y (nx502), .A0 (\output [8]), .A1 (\input [8]), .S0 (enable)
          ) ;
    dffr reg_output_9 (.Q (\output [9]), .QB (\$dummy [9]), .D (nx512), .CLK (
         clk), .R (nx845)) ;
    mux21 ix513 (.Y (nx512), .A0 (\output [9]), .A1 (\input [9]), .S0 (enable)
          ) ;
    dffr reg_output_10 (.Q (\output [10]), .QB (\$dummy [10]), .D (nx522), .CLK (
         clk), .R (nx845)) ;
    mux21 ix523 (.Y (nx522), .A0 (\output [10]), .A1 (\input [10]), .S0 (enable)
          ) ;
    dffr reg_output_11 (.Q (\output [11]), .QB (\$dummy [11]), .D (nx532), .CLK (
         clk), .R (nx845)) ;
    mux21 ix533 (.Y (nx532), .A0 (\output [11]), .A1 (\input [11]), .S0 (enable)
          ) ;
    dffr reg_output_12 (.Q (\output [12]), .QB (\$dummy [12]), .D (nx542), .CLK (
         clk), .R (nx845)) ;
    mux21 ix543 (.Y (nx542), .A0 (\output [12]), .A1 (\input [12]), .S0 (enable)
          ) ;
    dffr reg_output_13 (.Q (\output [13]), .QB (\$dummy [13]), .D (nx552), .CLK (
         clk), .R (nx845)) ;
    mux21 ix553 (.Y (nx552), .A0 (\output [13]), .A1 (\input [13]), .S0 (enable)
          ) ;
    dffr reg_output_14 (.Q (\output [14]), .QB (\$dummy [14]), .D (nx562), .CLK (
         clk), .R (nx845)) ;
    mux21 ix563 (.Y (nx562), .A0 (\output [14]), .A1 (\input [14]), .S0 (enable)
          ) ;
    dffr reg_output_15 (.Q (\output [15]), .QB (\$dummy [15]), .D (nx572), .CLK (
         clk), .R (nx847)) ;
    mux21 ix573 (.Y (nx572), .A0 (\output [15]), .A1 (\input [15]), .S0 (enable)
          ) ;
    dffr reg_output_16 (.Q (\output [16]), .QB (\$dummy [16]), .D (nx582), .CLK (
         clk), .R (nx847)) ;
    mux21 ix583 (.Y (nx582), .A0 (\output [16]), .A1 (\input [16]), .S0 (enable)
          ) ;
    dffr reg_output_17 (.Q (\output [17]), .QB (\$dummy [17]), .D (nx592), .CLK (
         clk), .R (nx847)) ;
    mux21 ix593 (.Y (nx592), .A0 (\output [17]), .A1 (\input [17]), .S0 (enable)
          ) ;
    dffr reg_output_18 (.Q (\output [18]), .QB (\$dummy [18]), .D (nx602), .CLK (
         clk), .R (nx847)) ;
    mux21 ix603 (.Y (nx602), .A0 (\output [18]), .A1 (\input [18]), .S0 (enable)
          ) ;
    dffr reg_output_19 (.Q (\output [19]), .QB (\$dummy [19]), .D (nx612), .CLK (
         clk), .R (nx847)) ;
    mux21 ix613 (.Y (nx612), .A0 (\output [19]), .A1 (\input [19]), .S0 (enable)
          ) ;
    dffr reg_output_20 (.Q (\output [20]), .QB (\$dummy [20]), .D (nx622), .CLK (
         clk), .R (nx847)) ;
    mux21 ix623 (.Y (nx622), .A0 (\output [20]), .A1 (\input [20]), .S0 (enable)
          ) ;
    dffr reg_output_21 (.Q (\output [21]), .QB (\$dummy [21]), .D (nx632), .CLK (
         clk), .R (nx847)) ;
    mux21 ix633 (.Y (nx632), .A0 (\output [21]), .A1 (\input [21]), .S0 (enable)
          ) ;
    dffr reg_output_22 (.Q (\output [22]), .QB (\$dummy [22]), .D (nx642), .CLK (
         clk), .R (nx847)) ;
    mux21 ix643 (.Y (nx642), .A0 (\output [22]), .A1 (\input [22]), .S0 (enable)
          ) ;
    dffr reg_output_23 (.Q (\output [23]), .QB (\$dummy [23]), .D (nx652), .CLK (
         clk), .R (nx847)) ;
    mux21 ix653 (.Y (nx652), .A0 (\output [23]), .A1 (\input [23]), .S0 (enable)
          ) ;
    dffr reg_output_24 (.Q (\output [24]), .QB (\$dummy [24]), .D (nx662), .CLK (
         clk), .R (nx847)) ;
    mux21 ix663 (.Y (nx662), .A0 (\output [24]), .A1 (\input [24]), .S0 (enable)
          ) ;
    dffr reg_output_25 (.Q (\output [25]), .QB (\$dummy [25]), .D (nx672), .CLK (
         clk), .R (nx847)) ;
    mux21 ix673 (.Y (nx672), .A0 (\output [25]), .A1 (\input [25]), .S0 (enable)
          ) ;
    dffr reg_output_26 (.Q (\output [26]), .QB (\$dummy [26]), .D (nx682), .CLK (
         clk), .R (nx847)) ;
    mux21 ix683 (.Y (nx682), .A0 (\output [26]), .A1 (\input [26]), .S0 (enable)
          ) ;
    dffr reg_output_27 (.Q (\output [27]), .QB (\$dummy [27]), .D (nx692), .CLK (
         clk), .R (nx847)) ;
    mux21 ix693 (.Y (nx692), .A0 (\output [27]), .A1 (\input [27]), .S0 (enable)
          ) ;
    dffr reg_output_28 (.Q (\output [28]), .QB (\$dummy [28]), .D (nx702), .CLK (
         clk), .R (nx847)) ;
    mux21 ix703 (.Y (nx702), .A0 (\output [28]), .A1 (\input [28]), .S0 (enable)
          ) ;
    dffr reg_output_29 (.Q (\output [29]), .QB (\$dummy [29]), .D (nx712), .CLK (
         clk), .R (nx847)) ;
    mux21 ix713 (.Y (nx712), .A0 (\output [29]), .A1 (\input [29]), .S0 (enable)
          ) ;
    dffr reg_output_30 (.Q (\output [30]), .QB (\$dummy [30]), .D (nx722), .CLK (
         clk), .R (NOT_reset)) ;
    mux21 ix723 (.Y (nx722), .A0 (\output [30]), .A1 (\input [30]), .S0 (enable)
          ) ;
    dffr reg_output_31 (.Q (\output [31]), .QB (\$dummy [31]), .D (nx732), .CLK (
         clk), .R (NOT_reset)) ;
    mux21 ix733 (.Y (nx732), .A0 (\output [31]), .A1 (\input [31]), .S0 (enable)
          ) ;
    inv01 ix844 (.Y (nx845), .A (reset)) ;
    inv01 ix846 (.Y (nx847), .A (reset)) ;
endmodule


module Multiplier_32 ( A, B, Product ) ;

    input [15:0]A ;
    input [15:0]B ;
    output [31:0]Product ;

    wire nx14, nx20, nx36, nx44, nx52, nx68, nx70, nx74, nx88, nx96, nx112, 
         nx114, nx122, nx128, nx144, nx152, nx168, nx170, nx180, nx188, nx196, 
         nx212, nx220, nx236, nx238, nx248, nx250, nx254, nx268, nx276, nx292, 
         nx300, nx316, nx318, nx328, nx330, nx338, nx344, nx360, nx368, nx384, 
         nx392, nx408, nx410, nx420, nx422, nx432, nx440, nx448, nx464, nx472, 
         nx488, nx496, nx512, nx514, nx524, nx526, nx536, nx538, nx542, nx556, 
         nx564, nx580, nx588, nx604, nx612, nx628, nx630, nx640, nx642, nx652, 
         nx654, nx662, nx668, nx684, nx692, nx708, nx716, nx732, nx740, nx756, 
         nx758, nx768, nx770, nx780, nx782, nx792, nx800, nx808, nx824, nx832, 
         nx848, nx856, nx872, nx880, nx896, nx898, nx908, nx910, nx920, nx922, 
         nx932, nx934, nx938, nx952, nx960, nx976, nx984, nx1000, nx1008, nx1024, 
         nx1032, nx1048, nx1050, nx1060, nx1062, nx1072, nx1074, nx1084, nx1086, 
         nx1094, nx1100, nx1116, nx1124, nx1140, nx1148, nx1164, nx1172, nx1188, 
         nx1196, nx1212, nx1214, nx1224, nx1226, nx1236, nx1238, nx1248, nx1250, 
         nx1260, nx1262, nx1268, nx1274, nx1290, nx1298, nx1314, nx1322, nx1338, 
         nx1346, nx1362, nx1370, nx1382, nx1390, nx1392, nx1402, nx1404, nx1414, 
         nx1416, nx1426, nx1428, nx1438, nx1440, nx1446, nx1452, nx1458, nx1466, 
         nx1474, nx1482, nx1490, nx1498, nx1506, nx1514, nx1522, nx1530, nx1538, 
         nx1546, nx1558, nx1560, nx1562, nx1564, nx1570, nx1572, nx1574, nx1576, 
         nx1582, nx1584, nx1586, nx1588, nx1594, nx1596, nx1598, nx1600, nx1602, 
         nx1604, nx1622, nx1630, nx1654, nx1662, nx1670, nx1678, nx1702, nx1710, 
         nx1718, nx1720, nx1734, nx1736, nx1738, nx1740, nx1742, nx1744, nx1758, 
         nx1760, nx1762, nx1764, nx1770, nx1776, nx1782, nx1790, nx1798, nx1830, 
         nx1838, nx1846, nx1854, nx1862, nx1870, nx1872, nx1874, nx1876, nx1882, 
         nx1884, nx1902, nx1904, nx1910, nx1912, nx1924, nx1938, nx1946, nx1954, 
         nx1962, nx1978, nx1986, nx1994, nx2002, nx2010, nx2012, nx2014, nx2016, 
         nx2018, nx2020, nx2030, nx2032, nx2038, nx2040, nx2048, nx2054, nx2060, 
         nx2074, nx2082, nx2090, nx2098, nx2106, nx2114, nx2122, nx2130, nx2138, 
         nx2140, nx2142, nx2144, nx2146, nx2148, nx2150, nx2152, nx2158, nx2160, 
         nx2162, nx2164, nx2170, nx2172, nx2184, nx2206, nx2214, nx2222, nx2230, 
         nx2238, nx2246, nx2254, nx2256, nx2258, nx2260, nx2262, nx2264, nx2266, 
         nx2268, nx2270, nx2272, nx2284, nx2290, nx2296, nx2302, nx2310, nx2318, 
         nx2326, nx2334, nx2342, nx2350, nx2358, nx2360, nx2362, nx2364, nx2366, 
         nx2368, nx2370, nx2372, nx2374, nx2376, nx2378, nx2380, nx2382, nx2384, 
         nx2402, nx2410, nx2418, nx2426, nx2434, nx2442, nx2450, nx2452, nx2454, 
         nx2456, nx2458, nx2460, nx2462, nx2464, nx2466, nx2468, nx2470, nx2472, 
         nx2478, nx2484, nx2490, nx2498, nx2506, nx2514, nx2522, nx2530, nx2532, 
         nx2534, nx2536, nx2538, nx2540, nx2542, nx2544, nx2546, nx2548, nx2566, 
         nx2574, nx2582, nx2590, nx2598, nx2600, nx2602, nx2604, nx2606, nx2608, 
         nx2610, nx2612, nx2618, nx2624, nx2630, nx2638, nx2646, nx2654, nx2656, 
         nx2658, nx2660, nx2662, nx2664, nx2682, nx2690, nx2698, nx2700, nx2702, 
         nx2704, nx2710, nx2716, nx2722, nx2730, nx2732, nx2738, nx2744, nx2748, 
         nx1551, nx1553, nx1559, nx1561, nx1563, nx1567, nx1569, nx1571, nx1573, 
         nx1579, nx1581, nx1583, nx1587, nx1589, nx1591, nx1593, nx1595, nx1597, 
         nx1599, nx1601, nx1605, nx1607, nx1611, nx1613, nx1615, nx1617, nx1621, 
         nx1627, nx1629, nx1631, nx1633, nx1635, nx1637, nx1639, nx1641, nx1643, 
         nx1645, nx1647, nx1653, nx1657, nx1659, nx1661, nx1667, nx1669, nx1671, 
         nx1673, nx1677, nx1679, nx1681, nx1683, nx1685, nx1687, nx1689, nx1691, 
         nx1693, nx1695, nx1699, nx1703, nx1709, nx1715, nx1717, nx1719, nx1721, 
         nx1723, nx1725, nx1727, nx1731, nx1733, nx1735, nx1737, nx1741, nx1743, 
         nx1749, nx1753, nx1755, nx1757, nx1763, nx1765, nx1767, nx1769, nx1773, 
         nx1775, nx1777, nx1779, nx1781, nx1785, nx1787, nx1789, nx1791, nx1795, 
         nx1799, nx1805, nx1807, nx1809, nx1811, nx1813, nx1815, nx1817, nx1821, 
         nx1825, nx1831, nx1837, nx1839, nx1841, nx1843, nx1845, nx1847, nx1849, 
         nx1851, nx1855, nx1857, nx1859, nx1865, nx1867, nx1871, nx1873, nx1879, 
         nx1883, nx1885, nx1887, nx1893, nx1895, nx1897, nx1899, nx1903, nx1905, 
         nx1907, nx1909, nx1911, nx1915, nx1917, nx1919, nx1921, nx1923, nx1927, 
         nx1933, nx1935, nx1937, nx1939, nx1941, nx1943, nx1945, nx1949, nx1953, 
         nx1959, nx1961, nx1963, nx1965, nx1967, nx1969, nx1971, nx1975, nx1979, 
         nx1985, nx1991, nx1993, nx1995, nx1997, nx1999, nx2001, nx2003, nx2005, 
         nx2011, nx2013, nx2017, nx2019, nx2025, nx2027, nx2031, nx2033, nx2039, 
         nx2043, nx2045, nx2047, nx2053, nx2055, nx2057, nx2059, nx2063, nx2065, 
         nx2067, nx2069, nx2071, nx2075, nx2077, nx2079, nx2081, nx2083, nx2087, 
         nx2089, nx2091, nx2093, nx2095, nx2097, nx2099, nx2101, nx2103, nx2105, 
         nx2109, nx2113, nx2119, nx2121, nx2123, nx2125, nx2127, nx2129, nx2131, 
         nx2135, nx2139, nx2145, nx2147, nx2149, nx2151, nx2153, nx2155, nx2157, 
         nx2161, nx2165, nx2171, nx2177, nx2179, nx2181, nx2183, nx2185, nx2187, 
         nx2189, nx2193, nx2195, nx2197, nx2199, nx2203, nx2205, nx2211, nx2213, 
         nx2217, nx2219, nx2225, nx2227, nx2231, nx2233, nx2239, nx2243, nx2245, 
         nx2247, nx2253, nx2255, nx2257, nx2259, nx2263, nx2265, nx2267, nx2269, 
         nx2271, nx2275, nx2277, nx2279, nx2281, nx2283, nx2287, nx2289, nx2291, 
         nx2293, nx2295, nx2299, nx2301, nx2303, nx2305, nx2309, nx2313, nx2319, 
         nx2321, nx2323, nx2325, nx2327, nx2329, nx2331, nx2335, nx2339, nx2345, 
         nx2347, nx2349, nx2351, nx2353, nx2355, nx2357, nx2361, nx2365, nx2371, 
         nx2373, nx2375, nx2377, nx2379, nx2381, nx2383, nx2387, nx2391, nx2397, 
         nx2403, nx2405, nx2407, nx2409, nx2411, nx2413, nx2415, nx2419, nx2423, 
         nx2427, nx2431, nx2435, nx2439, nx2443, nx2447, nx2451, nx2453, nx2455, 
         nx2461, nx2465, nx2469, nx2473, nx2479, nx2481, nx2483, nx2485, nx2487, 
         nx2489, nx2491, nx2493, nx2497, nx2501, nx2507, nx2509, nx2511, nx2513, 
         nx2515, nx2517, nx2519, nx2523, nx2527, nx2533, nx2535, nx2537, nx2539, 
         nx2541, nx2543, nx2545, nx2549, nx2553, nx2559, nx2561, nx2563, nx2565, 
         nx2567, nx2569, nx2571, nx2575, nx2579, nx2585, nx2591, nx2593, nx2595, 
         nx2597, nx2599, nx2601, nx2603, nx2607, nx2637, nx2639, nx2643, nx2645, 
         nx2651, nx2653, nx2655, nx2657, nx2659, nx2661, nx2663, nx2667, nx2671, 
         nx2677, nx2679, nx2681, nx2683, nx2685, nx2687, nx2689, nx2693, nx2697, 
         nx2703, nx2705, nx2707, nx2709, nx2711, nx2713, nx2715, nx2719, nx2723, 
         nx2729, nx2731, nx2733, nx2735, nx2737, nx2739, nx2741, nx2745, nx2749, 
         nx2755, nx2761, nx2763, nx2765, nx2767, nx2769, nx2775, nx2785, nx2787, 
         nx2793, nx2797, nx2801, nx2807, nx2809, nx2811, nx2813, nx2819, nx2823, 
         nx2827, nx2833, nx2835, nx2837, nx2839, nx2845, nx2849, nx2853, nx2859, 
         nx2861, nx2863, nx2865, nx2871, nx2875, nx2879, nx2883, nx2887, nx2889, 
         nx2891, nx2893, nx2895, nx2897, nx2900, nx2907, nx2910, nx2914, nx2918, 
         nx2920, nx2924, nx2926, nx2928, nx2930, nx2932, nx2934, nx2936, nx2938, 
         nx2941, nx2943, nx2945, nx2948, nx2950, nx2955, nx2958, nx2961, nx2964, 
         nx2968, nx2972, nx2974, nx2978, nx2980, nx2982, nx2984, nx2986, nx2988, 
         nx2990, nx2992, nx2995, nx2997, nx2999, nx3002, nx3004, nx3007, nx3011, 
         nx3015, nx3017, nx3019, nx3023, nx3025, nx3028, nx3033, nx3037, nx3039, 
         nx3041, nx3045, nx3049, nx3051, nx3053, nx3055, nx3057, nx3059, nx3061, 
         nx3063, nx3066, nx3068, nx3070, nx3072, nx3075, nx3077, nx3079, nx3082, 
         nx3087, nx3091, nx3093, nx3095, nx3099, nx3102, nx3105, nx3109, nx3111, 
         nx3113, nx3115, nx3118, nx3123, nx3127, nx3129, nx3131, nx3133, nx3135, 
         nx3138, nx3141, nx3145, nx3147, nx3149, nx3153, nx3157, nx3159, nx3161, 
         nx3163, nx3165, nx3167, nx3169, nx3172, nx3175, nx3178, nx3181, nx3184, 
         nx3188, nx3192, nx3196, nx3198, nx3200, nx3204, nx3206, nx3212, nx3214, 
         nx3216, nx3218, nx3220, nx3223, nx3226, nx3229, nx3232, nx3236, nx3238, 
         nx3240, nx3242, nx3246, nx3249, nx3252, nx3255, nx3259, nx3262, nx3266, 
         nx3270, nx3274, nx3276, nx3278, nx3281, nx3286, nx3288, nx3290, nx3292, 
         nx3294, nx3296, nx3299, nx3301, nx3303, nx3306, nx3311, nx3314, nx3317, 
         nx3320, nx3324, nx3327, nx3331, nx3334, nx3338, nx3342, nx3346, nx3348, 
         nx3350, nx3354, nx3356, nx3360, nx3364, nx3367, nx3370, nx3373, nx3377, 
         nx3380, nx3384, nx3387, nx3391, nx3394, nx3398, nx3402, nx3406, nx3408, 
         nx3410, nx3413, nx3417, nx3420, nx3424, nx3427, nx3431, nx3434, nx3438, 
         nx3441, nx3445, nx3448, nx3452, nx3456, nx3460, nx3462, nx3464, nx3468, 
         nx3470, nx3473, nx3477, nx3481, nx3484, nx3488, nx3491, nx3495, nx3498, 
         nx3502, nx3506, nx3510, nx3512, nx3514, nx3517, nx3521, nx3525, nx3529, 
         nx3532, nx3536, nx3539, nx3543, nx3547, nx3551, nx3553, nx3555, nx3559, 
         nx3561, nx3564, nx3568, nx3572, nx3575, nx3579, nx3583, nx3587, nx3589, 
         nx3591, nx3594, nx3598, nx3602, nx3606, nx3610, nx3614, nx3616, nx3618, 
         nx3622, nx3624, nx3627, nx3632, nx3636, nx3638, nx3640, nx3643, nx3648, 
         nx3652, nx3665, nx3667, nx3669, nx3671, nx3673, nx3675, nx3677, nx3679, 
         nx3681, nx3683, nx3685, nx3687, nx3689, nx3691, nx3693, nx3695, nx3697, 
         nx3699, nx3701, nx3703, nx3705, nx3707, nx3709, nx3711, nx3713, nx3715, 
         nx3717, nx3719, nx3721, nx3723, nx3725, nx3727, nx3729, nx3731, nx3733, 
         nx3735, nx3737, nx3739, nx3741, nx3743, nx3745, nx3747, nx3749, nx3751, 
         nx3753, nx3755, nx3757, nx3759, nx3761, nx3763, nx3765, nx3767, nx3769, 
         nx3771, nx3773, nx3775, nx3777, nx3779, nx3781, nx3783, nx3785, nx3787, 
         nx3789, nx3791;



    xor2 ix2791 (.Y (Product[15]), .A0 (nx1094), .A1 (nx1260)) ;
    nor02ii ix1095 (.Y (nx1094), .A0 (nx1551), .A1 (nx938)) ;
    xnor2 ix1552 (.Y (nx1551), .A0 (nx1553), .A1 (nx2301)) ;
    aoi32 ix1554 (.Y (nx1553), .A0 (nx3737), .A1 (nx3725), .A2 (nx932), .B0 (
          nx800), .B1 (nx934)) ;
    xnor2 ix933 (.Y (nx932), .A0 (nx808), .A1 (nx2093)) ;
    oai32 ix809 (.Y (nx808), .A0 (nx1559), .A1 (nx1561), .A2 (nx1563), .B0 (
          nx2005), .B1 (nx2089)) ;
    inv01 ix1560 (.Y (nx1559), .A (B[11])) ;
    inv01 ix1562 (.Y (nx1561), .A (A[1])) ;
    xnor2 ix1564 (.Y (nx1563), .A0 (nx684), .A1 (nx782)) ;
    oai32 ix685 (.Y (nx684), .A0 (nx1567), .A1 (nx1569), .A2 (nx1571), .B0 (
          nx1851), .B1 (nx1921)) ;
    inv01 ix1568 (.Y (nx1567), .A (B[9])) ;
    inv01 ix1570 (.Y (nx1569), .A (A[2])) ;
    xnor2 ix1572 (.Y (nx1571), .A0 (nx1573), .A1 (nx1787)) ;
    aoi32 ix1574 (.Y (nx1573), .A0 (nx3761), .A1 (nx3713), .A2 (nx524), .B0 (
          nx464), .B1 (nx526)) ;
    xnor2 ix525 (.Y (nx524), .A0 (nx472), .A1 (nx1683)) ;
    oai32 ix473 (.Y (nx472), .A0 (nx1579), .A1 (nx1581), .A2 (nx1583), .B0 (
          nx1647), .B1 (nx1679)) ;
    inv02 ix1580 (.Y (nx1579), .A (B[5])) ;
    inv02 ix1582 (.Y (nx1581), .A (A[4])) ;
    xnor2 ix1584 (.Y (nx1583), .A0 (nx384), .A1 (nx410)) ;
    oai32 ix385 (.Y (nx384), .A0 (nx1587), .A1 (nx1589), .A2 (nx1591), .B0 (
          nx1601), .B1 (nx1615)) ;
    inv02 ix1588 (.Y (nx1587), .A (B[3])) ;
    inv01 ix1590 (.Y (nx1589), .A (A[5])) ;
    xnor2 ix1592 (.Y (nx1591), .A0 (nx1593), .A1 (nx1595)) ;
    nand02 ix1594 (.Y (nx1593), .A0 (nx3781), .A1 (nx3701)) ;
    xnor2 ix1596 (.Y (nx1595), .A0 (nx1597), .A1 (nx1599)) ;
    nand02 ix1598 (.Y (nx1597), .A0 (nx3785), .A1 (nx3697)) ;
    nand02 ix1600 (.Y (nx1599), .A0 (nx3693), .A1 (nx3789)) ;
    inv01 ix1606 (.Y (nx1605), .A (A[7])) ;
    inv01 ix1608 (.Y (nx1607), .A (B[0])) ;
    nand02 ix1612 (.Y (nx1611), .A0 (nx3785), .A1 (nx3701)) ;
    nand02 ix1614 (.Y (nx1613), .A0 (nx3697), .A1 (nx3789)) ;
    xnor2 ix1616 (.Y (nx1615), .A0 (nx1617), .A1 (nx1591)) ;
    nand02 ix1618 (.Y (nx1617), .A0 (nx3777), .A1 (nx3705)) ;
    xnor2 ix411 (.Y (nx410), .A0 (nx1621), .A1 (nx408)) ;
    nand02 ix1622 (.Y (nx1621), .A0 (nx3773), .A1 (nx3705)) ;
    xnor2 ix409 (.Y (nx408), .A0 (nx392), .A1 (nx1633)) ;
    oai33 ix393 (.Y (nx392), .A0 (nx1627), .A1 (nx1629), .A2 (nx1595), .B0 (
          nx1631), .B1 (nx1605), .B2 (nx1599)) ;
    inv02 ix1628 (.Y (nx1627), .A (B[2])) ;
    inv01 ix1630 (.Y (nx1629), .A (A[6])) ;
    inv02 ix1632 (.Y (nx1631), .A (B[1])) ;
    xnor2 ix1634 (.Y (nx1633), .A0 (nx1635), .A1 (nx1637)) ;
    nand02 ix1636 (.Y (nx1635), .A0 (nx3777), .A1 (nx3701)) ;
    xnor2 ix1638 (.Y (nx1637), .A0 (nx1639), .A1 (nx1641)) ;
    nand02 ix1640 (.Y (nx1639), .A0 (nx3781), .A1 (nx3697)) ;
    xnor2 ix1642 (.Y (nx1641), .A0 (nx1643), .A1 (nx1645)) ;
    nand02 ix1644 (.Y (nx1643), .A0 (nx3785), .A1 (nx3693)) ;
    nand02 ix1646 (.Y (nx1645), .A0 (nx3689), .A1 (nx3789)) ;
    aoi32 ix1648 (.Y (nx1647), .A0 (nx3773), .A1 (nx3709), .A2 (nx316), .B0 (
          nx292), .B1 (nx318)) ;
    xnor2 ix317 (.Y (nx316), .A0 (nx300), .A1 (nx1615)) ;
    oai33 ix301 (.Y (nx300), .A0 (nx1627), .A1 (nx1589), .A2 (nx1653), .B0 (
          nx1631), .B1 (nx1629), .B2 (nx1613)) ;
    xnor2 ix1654 (.Y (nx1653), .A0 (nx1611), .A1 (nx1613)) ;
    oai32 ix293 (.Y (nx292), .A0 (nx1587), .A1 (nx1581), .A2 (nx1657), .B0 (
          nx1661), .B1 (nx1671)) ;
    xnor2 ix1658 (.Y (nx1657), .A0 (nx1659), .A1 (nx1653)) ;
    nand02 ix1660 (.Y (nx1659), .A0 (nx3781), .A1 (nx3705)) ;
    nand02 ix1668 (.Y (nx1667), .A0 (nx3785), .A1 (nx3705)) ;
    nand02 ix1670 (.Y (nx1669), .A0 (nx3701), .A1 (nx3789)) ;
    xnor2 ix1672 (.Y (nx1671), .A0 (nx1673), .A1 (nx1657)) ;
    nand02 ix1674 (.Y (nx1673), .A0 (nx3777), .A1 (nx3709)) ;
    xnor2 ix319 (.Y (nx318), .A0 (nx1677), .A1 (nx316)) ;
    nand02 ix1678 (.Y (nx1677), .A0 (nx3773), .A1 (nx3709)) ;
    xnor2 ix1680 (.Y (nx1679), .A0 (nx1681), .A1 (nx1583)) ;
    nand02 ix1682 (.Y (nx1681), .A0 (nx3769), .A1 (nx3709)) ;
    xnor2 ix1684 (.Y (nx1683), .A0 (nx1685), .A1 (nx1687)) ;
    nand02 ix1686 (.Y (nx1685), .A0 (nx3765), .A1 (nx3709)) ;
    xnor2 ix1688 (.Y (nx1687), .A0 (nx1689), .A1 (nx1691)) ;
    aoi32 ix1690 (.Y (nx1689), .A0 (nx3773), .A1 (nx3705), .A2 (nx408), .B0 (
          nx384), .B1 (nx410)) ;
    xnor2 ix1692 (.Y (nx1691), .A0 (nx1693), .A1 (nx1695)) ;
    nand02 ix1694 (.Y (nx1693), .A0 (nx3769), .A1 (nx3705)) ;
    xnor2 ix1696 (.Y (nx1695), .A0 (nx488), .A1 (nx514)) ;
    oai32 ix489 (.Y (nx488), .A0 (nx1587), .A1 (nx1629), .A2 (nx1637), .B0 (
          nx1699), .B1 (nx1633)) ;
    inv01 ix1704 (.Y (nx1703), .A (A[8])) ;
    xnor2 ix515 (.Y (nx514), .A0 (nx1709), .A1 (nx512)) ;
    nand02 ix1710 (.Y (nx1709), .A0 (nx3773), .A1 (nx3701)) ;
    xnor2 ix513 (.Y (nx512), .A0 (nx496), .A1 (nx1715)) ;
    oai33 ix497 (.Y (nx496), .A0 (nx1627), .A1 (nx1605), .A2 (nx1641), .B0 (
          nx1631), .B1 (nx1703), .B2 (nx1645)) ;
    xnor2 ix1716 (.Y (nx1715), .A0 (nx1717), .A1 (nx1719)) ;
    nand02 ix1718 (.Y (nx1717), .A0 (nx3777), .A1 (nx3697)) ;
    xnor2 ix1720 (.Y (nx1719), .A0 (nx1721), .A1 (nx1723)) ;
    nand02 ix1722 (.Y (nx1721), .A0 (nx3781), .A1 (nx3693)) ;
    xnor2 ix1724 (.Y (nx1723), .A0 (nx1725), .A1 (nx1727)) ;
    nand02 ix1726 (.Y (nx1725), .A0 (nx3785), .A1 (nx3689)) ;
    nand02 ix1728 (.Y (nx1727), .A0 (nx3685), .A1 (nx3789)) ;
    oai32 ix465 (.Y (nx464), .A0 (nx1731), .A1 (nx1733), .A2 (nx1735), .B0 (
          nx1737), .B1 (nx1779)) ;
    inv02 ix1732 (.Y (nx1731), .A (B[6])) ;
    inv01 ix1734 (.Y (nx1733), .A (A[3])) ;
    xnor2 ix1736 (.Y (nx1735), .A0 (nx1647), .A1 (nx1679)) ;
    inv01 ix1738 (.Y (nx1737), .A (nx368)) ;
    oai32 ix369 (.Y (nx368), .A0 (nx1579), .A1 (nx1733), .A2 (nx1741), .B0 (
          nx1743), .B1 (nx1775)) ;
    xnor2 ix1742 (.Y (nx1741), .A0 (nx292), .A1 (nx318)) ;
    aoi32 ix1744 (.Y (nx1743), .A0 (nx3773), .A1 (nx3713), .A2 (nx236), .B0 (
          nx212), .B1 (nx238)) ;
    xnor2 ix237 (.Y (nx236), .A0 (nx220), .A1 (nx1671)) ;
    oai33 ix221 (.Y (nx220), .A0 (nx1627), .A1 (nx1581), .A2 (nx1749), .B0 (
          nx1631), .B1 (nx1589), .B2 (nx1669)) ;
    xnor2 ix1750 (.Y (nx1749), .A0 (nx1667), .A1 (nx1669)) ;
    oai32 ix213 (.Y (nx212), .A0 (nx1587), .A1 (nx1733), .A2 (nx1753), .B0 (
          nx1757), .B1 (nx1767)) ;
    xnor2 ix1754 (.Y (nx1753), .A0 (nx1755), .A1 (nx1749)) ;
    nand02 ix1756 (.Y (nx1755), .A0 (nx3781), .A1 (nx3709)) ;
    nand02 ix1764 (.Y (nx1763), .A0 (nx3785), .A1 (nx3709)) ;
    nand02 ix1766 (.Y (nx1765), .A0 (nx3705), .A1 (nx3789)) ;
    xnor2 ix1768 (.Y (nx1767), .A0 (nx1769), .A1 (nx1753)) ;
    nand02 ix1770 (.Y (nx1769), .A0 (nx3777), .A1 (nx3713)) ;
    xnor2 ix239 (.Y (nx238), .A0 (nx1773), .A1 (nx236)) ;
    nand02 ix1774 (.Y (nx1773), .A0 (nx3773), .A1 (nx3713)) ;
    xnor2 ix1776 (.Y (nx1775), .A0 (nx1777), .A1 (nx1741)) ;
    nand02 ix1778 (.Y (nx1777), .A0 (nx3769), .A1 (nx3713)) ;
    xnor2 ix1780 (.Y (nx1779), .A0 (nx1781), .A1 (nx1735)) ;
    nand02 ix1782 (.Y (nx1781), .A0 (nx3765), .A1 (nx3713)) ;
    xnor2 ix527 (.Y (nx526), .A0 (nx1785), .A1 (nx524)) ;
    nand02 ix1786 (.Y (nx1785), .A0 (nx3761), .A1 (nx3713)) ;
    xnor2 ix1788 (.Y (nx1787), .A0 (nx1789), .A1 (nx1791)) ;
    nand02 ix1790 (.Y (nx1789), .A0 (nx3757), .A1 (nx3713)) ;
    xnor2 ix1792 (.Y (nx1791), .A0 (nx580), .A1 (nx642)) ;
    oai32 ix581 (.Y (nx580), .A0 (nx1731), .A1 (nx1581), .A2 (nx1687), .B0 (
          nx1795), .B1 (nx1683)) ;
    inv01 ix1796 (.Y (nx1795), .A (nx472)) ;
    xnor2 ix643 (.Y (nx642), .A0 (nx1799), .A1 (nx640)) ;
    nand02 ix1800 (.Y (nx1799), .A0 (nx3761), .A1 (nx3709)) ;
    xnor2 ix641 (.Y (nx640), .A0 (nx588), .A1 (nx1805)) ;
    oai32 ix589 (.Y (nx588), .A0 (nx1579), .A1 (nx1589), .A2 (nx1695), .B0 (
          nx1689), .B1 (nx1691)) ;
    xnor2 ix1806 (.Y (nx1805), .A0 (nx1807), .A1 (nx1809)) ;
    nand02 ix1808 (.Y (nx1807), .A0 (nx3765), .A1 (nx3705)) ;
    xnor2 ix1810 (.Y (nx1809), .A0 (nx1811), .A1 (nx1813)) ;
    aoi32 ix1812 (.Y (nx1811), .A0 (nx3773), .A1 (nx3701), .A2 (nx512), .B0 (
          nx488), .B1 (nx514)) ;
    xnor2 ix1814 (.Y (nx1813), .A0 (nx1815), .A1 (nx1817)) ;
    nand02 ix1816 (.Y (nx1815), .A0 (nx3769), .A1 (nx3701)) ;
    xnor2 ix1818 (.Y (nx1817), .A0 (nx604), .A1 (nx630)) ;
    oai32 ix605 (.Y (nx604), .A0 (nx1587), .A1 (nx1605), .A2 (nx1719), .B0 (
          nx1821), .B1 (nx1715)) ;
    inv01 ix1826 (.Y (nx1825), .A (A[9])) ;
    xnor2 ix631 (.Y (nx630), .A0 (nx1831), .A1 (nx628)) ;
    nand02 ix1832 (.Y (nx1831), .A0 (nx3773), .A1 (nx3697)) ;
    xnor2 ix629 (.Y (nx628), .A0 (nx612), .A1 (nx1837)) ;
    oai33 ix613 (.Y (nx612), .A0 (nx1627), .A1 (nx1703), .A2 (nx1723), .B0 (
          nx1631), .B1 (nx1825), .B2 (nx1727)) ;
    xnor2 ix1838 (.Y (nx1837), .A0 (nx1839), .A1 (nx1841)) ;
    nand02 ix1840 (.Y (nx1839), .A0 (nx3777), .A1 (nx3693)) ;
    xnor2 ix1842 (.Y (nx1841), .A0 (nx1843), .A1 (nx1845)) ;
    nand02 ix1844 (.Y (nx1843), .A0 (nx3781), .A1 (nx3689)) ;
    xnor2 ix1846 (.Y (nx1845), .A0 (nx1847), .A1 (nx1849)) ;
    nand02 ix1848 (.Y (nx1847), .A0 (nx3785), .A1 (nx3685)) ;
    nand02 ix1850 (.Y (nx1849), .A0 (nx3681), .A1 (nx3789)) ;
    inv01 ix1852 (.Y (nx1851), .A (nx564)) ;
    oai32 ix565 (.Y (nx564), .A0 (nx1855), .A1 (nx1569), .A2 (nx1857), .B0 (
          nx1859), .B1 (nx1917)) ;
    inv01 ix1856 (.Y (nx1855), .A (B[8])) ;
    xnor2 ix1858 (.Y (nx1857), .A0 (nx464), .A1 (nx526)) ;
    aoi32 ix1860 (.Y (nx1859), .A0 (nx3761), .A1 (nx3717), .A2 (nx420), .B0 (
          nx360), .B1 (nx422)) ;
    xnor2 ix421 (.Y (nx420), .A0 (nx368), .A1 (nx1779)) ;
    oai32 ix361 (.Y (nx360), .A0 (nx1731), .A1 (nx1569), .A2 (nx1865), .B0 (
          nx1867), .B1 (nx1909)) ;
    xnor2 ix1866 (.Y (nx1865), .A0 (nx1743), .A1 (nx1775)) ;
    inv01 ix1868 (.Y (nx1867), .A (nx276)) ;
    oai32 ix277 (.Y (nx276), .A0 (nx1579), .A1 (nx1569), .A2 (nx1871), .B0 (
          nx1873), .B1 (nx1905)) ;
    xnor2 ix1872 (.Y (nx1871), .A0 (nx212), .A1 (nx238)) ;
    aoi32 ix1874 (.Y (nx1873), .A0 (nx3773), .A1 (nx3717), .A2 (nx168), .B0 (
          nx144), .B1 (nx170)) ;
    xnor2 ix169 (.Y (nx168), .A0 (nx152), .A1 (nx1767)) ;
    oai33 ix153 (.Y (nx152), .A0 (nx1627), .A1 (nx1733), .A2 (nx1879), .B0 (
          nx1631), .B1 (nx1581), .B2 (nx1765)) ;
    xnor2 ix1880 (.Y (nx1879), .A0 (nx1763), .A1 (nx1765)) ;
    oai32 ix145 (.Y (nx144), .A0 (nx1587), .A1 (nx1569), .A2 (nx1883), .B0 (
          nx1887), .B1 (nx1897)) ;
    xnor2 ix1884 (.Y (nx1883), .A0 (nx1885), .A1 (nx1879)) ;
    nand02 ix1886 (.Y (nx1885), .A0 (nx3781), .A1 (nx3713)) ;
    nand02 ix1894 (.Y (nx1893), .A0 (nx3785), .A1 (nx3713)) ;
    nand02 ix1896 (.Y (nx1895), .A0 (nx3709), .A1 (nx3789)) ;
    xnor2 ix1898 (.Y (nx1897), .A0 (nx1899), .A1 (nx1883)) ;
    nand02 ix1900 (.Y (nx1899), .A0 (nx3777), .A1 (nx3717)) ;
    xnor2 ix171 (.Y (nx170), .A0 (nx1903), .A1 (nx168)) ;
    nand02 ix1904 (.Y (nx1903), .A0 (nx3773), .A1 (nx3717)) ;
    xnor2 ix1906 (.Y (nx1905), .A0 (nx1907), .A1 (nx1871)) ;
    nand02 ix1908 (.Y (nx1907), .A0 (nx3769), .A1 (nx3717)) ;
    xnor2 ix1910 (.Y (nx1909), .A0 (nx1911), .A1 (nx1865)) ;
    nand02 ix1912 (.Y (nx1911), .A0 (nx3765), .A1 (nx3717)) ;
    xnor2 ix423 (.Y (nx422), .A0 (nx1915), .A1 (nx420)) ;
    nand02 ix1916 (.Y (nx1915), .A0 (nx3761), .A1 (nx3717)) ;
    xnor2 ix1918 (.Y (nx1917), .A0 (nx1919), .A1 (nx1857)) ;
    nand02 ix1920 (.Y (nx1919), .A0 (nx3757), .A1 (nx3717)) ;
    xnor2 ix1922 (.Y (nx1921), .A0 (nx1923), .A1 (nx1571)) ;
    nand02 ix1924 (.Y (nx1923), .A0 (nx3753), .A1 (nx3717)) ;
    xnor2 ix783 (.Y (nx782), .A0 (nx1927), .A1 (nx780)) ;
    nand02 ix1928 (.Y (nx1927), .A0 (nx3749), .A1 (nx3717)) ;
    xnor2 ix781 (.Y (nx780), .A0 (nx692), .A1 (nx1933)) ;
    oai32 ix693 (.Y (nx692), .A0 (nx1855), .A1 (nx1733), .A2 (nx1791), .B0 (
          nx1573), .B1 (nx1787)) ;
    xnor2 ix1934 (.Y (nx1933), .A0 (nx1935), .A1 (nx1937)) ;
    nand02 ix1936 (.Y (nx1935), .A0 (nx3753), .A1 (nx3713)) ;
    xnor2 ix1938 (.Y (nx1937), .A0 (nx1939), .A1 (nx1941)) ;
    aoi32 ix1940 (.Y (nx1939), .A0 (nx3761), .A1 (nx3709), .A2 (nx640), .B0 (
          nx580), .B1 (nx642)) ;
    xnor2 ix1942 (.Y (nx1941), .A0 (nx1943), .A1 (nx1945)) ;
    nand02 ix1944 (.Y (nx1943), .A0 (nx3757), .A1 (nx3709)) ;
    xnor2 ix1946 (.Y (nx1945), .A0 (nx708), .A1 (nx770)) ;
    oai32 ix709 (.Y (nx708), .A0 (nx1731), .A1 (nx1589), .A2 (nx1809), .B0 (
          nx1949), .B1 (nx1805)) ;
    inv01 ix1950 (.Y (nx1949), .A (nx588)) ;
    xnor2 ix771 (.Y (nx770), .A0 (nx1953), .A1 (nx768)) ;
    nand02 ix1954 (.Y (nx1953), .A0 (nx3761), .A1 (nx3705)) ;
    xnor2 ix769 (.Y (nx768), .A0 (nx716), .A1 (nx1959)) ;
    oai32 ix717 (.Y (nx716), .A0 (nx1579), .A1 (nx1629), .A2 (nx1817), .B0 (
          nx1811), .B1 (nx1813)) ;
    xnor2 ix1960 (.Y (nx1959), .A0 (nx1961), .A1 (nx1963)) ;
    nand02 ix1962 (.Y (nx1961), .A0 (nx3765), .A1 (nx3701)) ;
    xnor2 ix1964 (.Y (nx1963), .A0 (nx1965), .A1 (nx1967)) ;
    aoi32 ix1966 (.Y (nx1965), .A0 (nx3773), .A1 (nx3697), .A2 (nx628), .B0 (
          nx604), .B1 (nx630)) ;
    xnor2 ix1968 (.Y (nx1967), .A0 (nx1969), .A1 (nx1971)) ;
    nand02 ix1970 (.Y (nx1969), .A0 (nx3769), .A1 (nx3697)) ;
    xnor2 ix1972 (.Y (nx1971), .A0 (nx732), .A1 (nx758)) ;
    oai32 ix733 (.Y (nx732), .A0 (nx1587), .A1 (nx1703), .A2 (nx1841), .B0 (
          nx1975), .B1 (nx1837)) ;
    inv01 ix1980 (.Y (nx1979), .A (A[10])) ;
    xnor2 ix759 (.Y (nx758), .A0 (nx1985), .A1 (nx756)) ;
    nand02 ix1986 (.Y (nx1985), .A0 (nx3773), .A1 (nx3693)) ;
    xnor2 ix757 (.Y (nx756), .A0 (nx740), .A1 (nx1991)) ;
    oai33 ix741 (.Y (nx740), .A0 (nx1627), .A1 (nx1825), .A2 (nx1845), .B0 (
          nx1631), .B1 (nx1979), .B2 (nx1849)) ;
    xnor2 ix1992 (.Y (nx1991), .A0 (nx1993), .A1 (nx1995)) ;
    nand02 ix1994 (.Y (nx1993), .A0 (nx3777), .A1 (nx3689)) ;
    xnor2 ix1996 (.Y (nx1995), .A0 (nx1997), .A1 (nx1999)) ;
    nand02 ix1998 (.Y (nx1997), .A0 (nx3781), .A1 (nx3685)) ;
    xnor2 ix2000 (.Y (nx1999), .A0 (nx2001), .A1 (nx2003)) ;
    nand02 ix2002 (.Y (nx2001), .A0 (nx3785), .A1 (nx3681)) ;
    nand02 ix2004 (.Y (nx2003), .A0 (nx3677), .A1 (nx3789)) ;
    aoi32 ix2006 (.Y (nx2005), .A0 (nx3749), .A1 (nx3721), .A2 (nx652), .B0 (
          nx556), .B1 (nx654)) ;
    xnor2 ix653 (.Y (nx652), .A0 (nx564), .A1 (nx1921)) ;
    oai32 ix557 (.Y (nx556), .A0 (nx1567), .A1 (nx1561), .A2 (nx2011), .B0 (
          nx2013), .B1 (nx2081)) ;
    xnor2 ix2012 (.Y (nx2011), .A0 (nx1859), .A1 (nx1917)) ;
    inv01 ix2014 (.Y (nx2013), .A (nx448)) ;
    oai32 ix449 (.Y (nx448), .A0 (nx1855), .A1 (nx1561), .A2 (nx2017), .B0 (
          nx2019), .B1 (nx2077)) ;
    xnor2 ix2018 (.Y (nx2017), .A0 (nx360), .A1 (nx422)) ;
    aoi32 ix2020 (.Y (nx2019), .A0 (nx3761), .A1 (nx3721), .A2 (nx328), .B0 (
          nx268), .B1 (nx330)) ;
    xnor2 ix329 (.Y (nx328), .A0 (nx276), .A1 (nx1909)) ;
    oai32 ix269 (.Y (nx268), .A0 (nx1731), .A1 (nx1561), .A2 (nx2025), .B0 (
          nx2027), .B1 (nx2069)) ;
    xnor2 ix2026 (.Y (nx2025), .A0 (nx1873), .A1 (nx1905)) ;
    inv01 ix2028 (.Y (nx2027), .A (nx196)) ;
    oai32 ix197 (.Y (nx196), .A0 (nx1579), .A1 (nx1561), .A2 (nx2031), .B0 (
          nx2033), .B1 (nx2065)) ;
    xnor2 ix2032 (.Y (nx2031), .A0 (nx144), .A1 (nx170)) ;
    aoi32 ix2034 (.Y (nx2033), .A0 (nx3773), .A1 (nx3721), .A2 (nx112), .B0 (
          nx88), .B1 (nx114)) ;
    xnor2 ix113 (.Y (nx112), .A0 (nx96), .A1 (nx1897)) ;
    oai33 ix97 (.Y (nx96), .A0 (nx1627), .A1 (nx1569), .A2 (nx2039), .B0 (nx1631
          ), .B1 (nx1733), .B2 (nx1895)) ;
    xnor2 ix2040 (.Y (nx2039), .A0 (nx1893), .A1 (nx1895)) ;
    oai32 ix89 (.Y (nx88), .A0 (nx1587), .A1 (nx1561), .A2 (nx2043), .B0 (nx2047
          ), .B1 (nx2057)) ;
    xnor2 ix2044 (.Y (nx2043), .A0 (nx2045), .A1 (nx2039)) ;
    nand02 ix2046 (.Y (nx2045), .A0 (nx3781), .A1 (nx3717)) ;
    nand02 ix2054 (.Y (nx2053), .A0 (nx3785), .A1 (nx3717)) ;
    nand02 ix2056 (.Y (nx2055), .A0 (nx3713), .A1 (nx3789)) ;
    xnor2 ix2058 (.Y (nx2057), .A0 (nx2059), .A1 (nx2043)) ;
    nand02 ix2060 (.Y (nx2059), .A0 (nx3777), .A1 (nx3721)) ;
    xnor2 ix115 (.Y (nx114), .A0 (nx2063), .A1 (nx112)) ;
    nand02 ix2064 (.Y (nx2063), .A0 (nx3773), .A1 (nx3721)) ;
    xnor2 ix2066 (.Y (nx2065), .A0 (nx2067), .A1 (nx2031)) ;
    nand02 ix2068 (.Y (nx2067), .A0 (nx3769), .A1 (nx3721)) ;
    xnor2 ix2070 (.Y (nx2069), .A0 (nx2071), .A1 (nx2025)) ;
    nand02 ix2072 (.Y (nx2071), .A0 (nx3765), .A1 (nx3721)) ;
    xnor2 ix331 (.Y (nx330), .A0 (nx2075), .A1 (nx328)) ;
    nand02 ix2076 (.Y (nx2075), .A0 (nx3761), .A1 (nx3721)) ;
    xnor2 ix2078 (.Y (nx2077), .A0 (nx2079), .A1 (nx2017)) ;
    nand02 ix2080 (.Y (nx2079), .A0 (nx3757), .A1 (nx3721)) ;
    xnor2 ix2082 (.Y (nx2081), .A0 (nx2083), .A1 (nx2011)) ;
    nand02 ix2084 (.Y (nx2083), .A0 (nx3753), .A1 (nx3721)) ;
    xnor2 ix655 (.Y (nx654), .A0 (nx2087), .A1 (nx652)) ;
    nand02 ix2088 (.Y (nx2087), .A0 (nx3749), .A1 (nx3721)) ;
    xnor2 ix2090 (.Y (nx2089), .A0 (nx2091), .A1 (nx1563)) ;
    nand02 ix2092 (.Y (nx2091), .A0 (nx3745), .A1 (nx3721)) ;
    xnor2 ix2094 (.Y (nx2093), .A0 (nx2095), .A1 (nx2097)) ;
    nand02 ix2096 (.Y (nx2095), .A0 (nx3741), .A1 (nx3721)) ;
    xnor2 ix2098 (.Y (nx2097), .A0 (nx2099), .A1 (nx2101)) ;
    aoi32 ix2100 (.Y (nx2099), .A0 (nx3749), .A1 (nx3717), .A2 (nx780), .B0 (
          nx684), .B1 (nx782)) ;
    xnor2 ix2102 (.Y (nx2101), .A0 (nx2103), .A1 (nx2105)) ;
    nand02 ix2104 (.Y (nx2103), .A0 (nx3745), .A1 (nx3717)) ;
    xnor2 ix2106 (.Y (nx2105), .A0 (nx824), .A1 (nx922)) ;
    oai32 ix825 (.Y (nx824), .A0 (nx1567), .A1 (nx1733), .A2 (nx1937), .B0 (
          nx2109), .B1 (nx1933)) ;
    inv01 ix2110 (.Y (nx2109), .A (nx692)) ;
    xnor2 ix923 (.Y (nx922), .A0 (nx2113), .A1 (nx920)) ;
    nand02 ix2114 (.Y (nx2113), .A0 (nx3749), .A1 (nx3713)) ;
    xnor2 ix921 (.Y (nx920), .A0 (nx832), .A1 (nx2119)) ;
    oai32 ix833 (.Y (nx832), .A0 (nx1855), .A1 (nx1581), .A2 (nx1945), .B0 (
          nx1939), .B1 (nx1941)) ;
    xnor2 ix2120 (.Y (nx2119), .A0 (nx2121), .A1 (nx2123)) ;
    nand02 ix2122 (.Y (nx2121), .A0 (nx3753), .A1 (nx3709)) ;
    xnor2 ix2124 (.Y (nx2123), .A0 (nx2125), .A1 (nx2127)) ;
    aoi32 ix2126 (.Y (nx2125), .A0 (nx3761), .A1 (nx3705), .A2 (nx768), .B0 (
          nx708), .B1 (nx770)) ;
    xnor2 ix2128 (.Y (nx2127), .A0 (nx2129), .A1 (nx2131)) ;
    nand02 ix2130 (.Y (nx2129), .A0 (nx3757), .A1 (nx3705)) ;
    xnor2 ix2132 (.Y (nx2131), .A0 (nx848), .A1 (nx910)) ;
    oai32 ix849 (.Y (nx848), .A0 (nx1731), .A1 (nx1629), .A2 (nx1963), .B0 (
          nx2135), .B1 (nx1959)) ;
    inv01 ix2136 (.Y (nx2135), .A (nx716)) ;
    xnor2 ix911 (.Y (nx910), .A0 (nx2139), .A1 (nx908)) ;
    nand02 ix2140 (.Y (nx2139), .A0 (nx3761), .A1 (nx3701)) ;
    xnor2 ix909 (.Y (nx908), .A0 (nx856), .A1 (nx2145)) ;
    oai32 ix857 (.Y (nx856), .A0 (nx1579), .A1 (nx1605), .A2 (nx1971), .B0 (
          nx1965), .B1 (nx1967)) ;
    xnor2 ix2146 (.Y (nx2145), .A0 (nx2147), .A1 (nx2149)) ;
    nand02 ix2148 (.Y (nx2147), .A0 (nx3765), .A1 (nx3697)) ;
    xnor2 ix2150 (.Y (nx2149), .A0 (nx2151), .A1 (nx2153)) ;
    aoi32 ix2152 (.Y (nx2151), .A0 (nx3775), .A1 (nx3693), .A2 (nx756), .B0 (
          nx732), .B1 (nx758)) ;
    xnor2 ix2154 (.Y (nx2153), .A0 (nx2155), .A1 (nx2157)) ;
    nand02 ix2156 (.Y (nx2155), .A0 (nx3769), .A1 (nx3693)) ;
    xnor2 ix2158 (.Y (nx2157), .A0 (nx872), .A1 (nx898)) ;
    oai32 ix873 (.Y (nx872), .A0 (nx1587), .A1 (nx1825), .A2 (nx1995), .B0 (
          nx2161), .B1 (nx1991)) ;
    inv01 ix2166 (.Y (nx2165), .A (A[11])) ;
    xnor2 ix899 (.Y (nx898), .A0 (nx2171), .A1 (nx896)) ;
    nand02 ix2172 (.Y (nx2171), .A0 (nx3775), .A1 (nx3689)) ;
    xnor2 ix897 (.Y (nx896), .A0 (nx880), .A1 (nx2177)) ;
    oai33 ix881 (.Y (nx880), .A0 (nx1627), .A1 (nx1979), .A2 (nx1999), .B0 (
          nx1631), .B1 (nx2165), .B2 (nx2003)) ;
    xnor2 ix2178 (.Y (nx2177), .A0 (nx2179), .A1 (nx2181)) ;
    nand02 ix2180 (.Y (nx2179), .A0 (nx3777), .A1 (nx3685)) ;
    xnor2 ix2182 (.Y (nx2181), .A0 (nx2183), .A1 (nx2185)) ;
    nand02 ix2184 (.Y (nx2183), .A0 (nx3781), .A1 (nx3681)) ;
    xnor2 ix2186 (.Y (nx2185), .A0 (nx2187), .A1 (nx2189)) ;
    nand02 ix2188 (.Y (nx2187), .A0 (nx3785), .A1 (nx3677)) ;
    nand02 ix2190 (.Y (nx2189), .A0 (nx3673), .A1 (nx3789)) ;
    oai32 ix801 (.Y (nx800), .A0 (nx2193), .A1 (nx2195), .A2 (nx2197), .B0 (
          nx2199), .B1 (nx2293)) ;
    inv01 ix2194 (.Y (nx2193), .A (B[12])) ;
    inv01 ix2196 (.Y (nx2195), .A (A[0])) ;
    xnor2 ix2198 (.Y (nx2197), .A0 (nx2005), .A1 (nx2089)) ;
    inv01 ix2200 (.Y (nx2199), .A (nx668)) ;
    oai32 ix669 (.Y (nx668), .A0 (nx1559), .A1 (nx2195), .A2 (nx2203), .B0 (
          nx2205), .B1 (nx2289)) ;
    xnor2 ix2204 (.Y (nx2203), .A0 (nx556), .A1 (nx654)) ;
    aoi32 ix2206 (.Y (nx2205), .A0 (nx3749), .A1 (nx3725), .A2 (nx536), .B0 (
          nx440), .B1 (nx538)) ;
    xnor2 ix537 (.Y (nx536), .A0 (nx448), .A1 (nx2081)) ;
    oai32 ix441 (.Y (nx440), .A0 (nx1567), .A1 (nx2195), .A2 (nx2211), .B0 (
          nx2213), .B1 (nx2281)) ;
    xnor2 ix2212 (.Y (nx2211), .A0 (nx2019), .A1 (nx2077)) ;
    inv01 ix2214 (.Y (nx2213), .A (nx344)) ;
    oai32 ix345 (.Y (nx344), .A0 (nx1855), .A1 (nx2195), .A2 (nx2217), .B0 (
          nx2219), .B1 (nx2277)) ;
    xnor2 ix2218 (.Y (nx2217), .A0 (nx268), .A1 (nx330)) ;
    aoi32 ix2220 (.Y (nx2219), .A0 (nx3761), .A1 (nx3725), .A2 (nx248), .B0 (
          nx188), .B1 (nx250)) ;
    xnor2 ix249 (.Y (nx248), .A0 (nx196), .A1 (nx2069)) ;
    oai32 ix189 (.Y (nx188), .A0 (nx1731), .A1 (nx2195), .A2 (nx2225), .B0 (
          nx2227), .B1 (nx2269)) ;
    xnor2 ix2226 (.Y (nx2225), .A0 (nx2033), .A1 (nx2065)) ;
    inv01 ix2228 (.Y (nx2227), .A (nx128)) ;
    oai32 ix129 (.Y (nx128), .A0 (nx1579), .A1 (nx2195), .A2 (nx2231), .B0 (
          nx2233), .B1 (nx2265)) ;
    xnor2 ix2232 (.Y (nx2231), .A0 (nx88), .A1 (nx114)) ;
    aoi32 ix2234 (.Y (nx2233), .A0 (nx3775), .A1 (nx3725), .A2 (nx68), .B0 (nx44
          ), .B1 (nx70)) ;
    xnor2 ix69 (.Y (nx68), .A0 (nx52), .A1 (nx2057)) ;
    oai33 ix53 (.Y (nx52), .A0 (nx1627), .A1 (nx1561), .A2 (nx2239), .B0 (nx1631
          ), .B1 (nx1569), .B2 (nx2055)) ;
    xnor2 ix2240 (.Y (nx2239), .A0 (nx2053), .A1 (nx2055)) ;
    oai32 ix45 (.Y (nx44), .A0 (nx1587), .A1 (nx2195), .A2 (nx2243), .B0 (nx2247
          ), .B1 (nx2257)) ;
    xnor2 ix2244 (.Y (nx2243), .A0 (nx2245), .A1 (nx2239)) ;
    nand02 ix2246 (.Y (nx2245), .A0 (nx3781), .A1 (nx3721)) ;
    nand02 ix2254 (.Y (nx2253), .A0 (nx3785), .A1 (nx3721)) ;
    nand02 ix2256 (.Y (nx2255), .A0 (nx3717), .A1 (nx3789)) ;
    xnor2 ix2258 (.Y (nx2257), .A0 (nx2259), .A1 (nx2243)) ;
    nand02 ix2260 (.Y (nx2259), .A0 (nx3777), .A1 (nx3725)) ;
    xnor2 ix71 (.Y (nx70), .A0 (nx2263), .A1 (nx68)) ;
    nand02 ix2264 (.Y (nx2263), .A0 (nx3775), .A1 (nx3725)) ;
    xnor2 ix2266 (.Y (nx2265), .A0 (nx2267), .A1 (nx2231)) ;
    nand02 ix2268 (.Y (nx2267), .A0 (nx3769), .A1 (nx3725)) ;
    xnor2 ix2270 (.Y (nx2269), .A0 (nx2271), .A1 (nx2225)) ;
    nand02 ix2272 (.Y (nx2271), .A0 (nx3765), .A1 (nx3725)) ;
    xnor2 ix251 (.Y (nx250), .A0 (nx2275), .A1 (nx248)) ;
    nand02 ix2276 (.Y (nx2275), .A0 (nx3761), .A1 (nx3725)) ;
    xnor2 ix2278 (.Y (nx2277), .A0 (nx2279), .A1 (nx2217)) ;
    nand02 ix2280 (.Y (nx2279), .A0 (nx3757), .A1 (nx3725)) ;
    xnor2 ix2282 (.Y (nx2281), .A0 (nx2283), .A1 (nx2211)) ;
    nand02 ix2284 (.Y (nx2283), .A0 (nx3753), .A1 (nx3725)) ;
    xnor2 ix539 (.Y (nx538), .A0 (nx2287), .A1 (nx536)) ;
    nand02 ix2288 (.Y (nx2287), .A0 (nx3749), .A1 (nx3725)) ;
    xnor2 ix2290 (.Y (nx2289), .A0 (nx2291), .A1 (nx2203)) ;
    nand02 ix2292 (.Y (nx2291), .A0 (nx3745), .A1 (nx3725)) ;
    xnor2 ix2294 (.Y (nx2293), .A0 (nx2295), .A1 (nx2197)) ;
    nand02 ix2296 (.Y (nx2295), .A0 (nx3741), .A1 (nx3725)) ;
    xnor2 ix935 (.Y (nx934), .A0 (nx2299), .A1 (nx932)) ;
    nand02 ix2300 (.Y (nx2299), .A0 (nx3737), .A1 (nx3725)) ;
    xnor2 ix2302 (.Y (nx2301), .A0 (nx2303), .A1 (nx2305)) ;
    nand02 ix2304 (.Y (nx2303), .A0 (nx3733), .A1 (nx3727)) ;
    xnor2 ix2306 (.Y (nx2305), .A0 (nx952), .A1 (nx1086)) ;
    oai32 ix953 (.Y (nx952), .A0 (nx2193), .A1 (nx1561), .A2 (nx2097), .B0 (
          nx2309), .B1 (nx2093)) ;
    inv01 ix2310 (.Y (nx2309), .A (nx808)) ;
    xnor2 ix1087 (.Y (nx1086), .A0 (nx2313), .A1 (nx1084)) ;
    nand02 ix2314 (.Y (nx2313), .A0 (nx3737), .A1 (nx3723)) ;
    xnor2 ix1085 (.Y (nx1084), .A0 (nx960), .A1 (nx2319)) ;
    oai32 ix961 (.Y (nx960), .A0 (nx1559), .A1 (nx1569), .A2 (nx2105), .B0 (
          nx2099), .B1 (nx2101)) ;
    xnor2 ix2320 (.Y (nx2319), .A0 (nx2321), .A1 (nx2323)) ;
    nand02 ix2322 (.Y (nx2321), .A0 (nx3741), .A1 (nx3719)) ;
    xnor2 ix2324 (.Y (nx2323), .A0 (nx2325), .A1 (nx2327)) ;
    aoi32 ix2326 (.Y (nx2325), .A0 (nx3749), .A1 (nx3713), .A2 (nx920), .B0 (
          nx824), .B1 (nx922)) ;
    xnor2 ix2328 (.Y (nx2327), .A0 (nx2329), .A1 (nx2331)) ;
    nand02 ix2330 (.Y (nx2329), .A0 (nx3745), .A1 (nx3713)) ;
    xnor2 ix2332 (.Y (nx2331), .A0 (nx976), .A1 (nx1074)) ;
    oai32 ix977 (.Y (nx976), .A0 (nx1567), .A1 (nx1581), .A2 (nx2123), .B0 (
          nx2335), .B1 (nx2119)) ;
    inv01 ix2336 (.Y (nx2335), .A (nx832)) ;
    xnor2 ix1075 (.Y (nx1074), .A0 (nx2339), .A1 (nx1072)) ;
    nand02 ix2340 (.Y (nx2339), .A0 (nx3749), .A1 (nx3709)) ;
    xnor2 ix1073 (.Y (nx1072), .A0 (nx984), .A1 (nx2345)) ;
    oai32 ix985 (.Y (nx984), .A0 (nx1855), .A1 (nx1589), .A2 (nx2131), .B0 (
          nx2125), .B1 (nx2127)) ;
    xnor2 ix2346 (.Y (nx2345), .A0 (nx2347), .A1 (nx2349)) ;
    nand02 ix2348 (.Y (nx2347), .A0 (nx3753), .A1 (nx3705)) ;
    xnor2 ix2350 (.Y (nx2349), .A0 (nx2351), .A1 (nx2353)) ;
    aoi32 ix2352 (.Y (nx2351), .A0 (nx3761), .A1 (nx3701), .A2 (nx908), .B0 (
          nx848), .B1 (nx910)) ;
    xnor2 ix2354 (.Y (nx2353), .A0 (nx2355), .A1 (nx2357)) ;
    nand02 ix2356 (.Y (nx2355), .A0 (nx3757), .A1 (nx3701)) ;
    xnor2 ix2358 (.Y (nx2357), .A0 (nx1000), .A1 (nx1062)) ;
    oai32 ix1001 (.Y (nx1000), .A0 (nx1731), .A1 (nx1605), .A2 (nx2149), .B0 (
          nx2361), .B1 (nx2145)) ;
    inv01 ix2362 (.Y (nx2361), .A (nx856)) ;
    xnor2 ix1063 (.Y (nx1062), .A0 (nx2365), .A1 (nx1060)) ;
    nand02 ix2366 (.Y (nx2365), .A0 (nx3761), .A1 (nx3697)) ;
    xnor2 ix1061 (.Y (nx1060), .A0 (nx1008), .A1 (nx2371)) ;
    oai32 ix1009 (.Y (nx1008), .A0 (nx1579), .A1 (nx1703), .A2 (nx2157), .B0 (
          nx2151), .B1 (nx2153)) ;
    xnor2 ix2372 (.Y (nx2371), .A0 (nx2373), .A1 (nx2375)) ;
    nand02 ix2374 (.Y (nx2373), .A0 (nx3765), .A1 (nx3693)) ;
    xnor2 ix2376 (.Y (nx2375), .A0 (nx2377), .A1 (nx2379)) ;
    aoi32 ix2378 (.Y (nx2377), .A0 (nx3775), .A1 (nx3689), .A2 (nx896), .B0 (
          nx872), .B1 (nx898)) ;
    xnor2 ix2380 (.Y (nx2379), .A0 (nx2381), .A1 (nx2383)) ;
    nand02 ix2382 (.Y (nx2381), .A0 (nx3769), .A1 (nx3689)) ;
    xnor2 ix2384 (.Y (nx2383), .A0 (nx1024), .A1 (nx1050)) ;
    oai32 ix1025 (.Y (nx1024), .A0 (nx1587), .A1 (nx1979), .A2 (nx2181), .B0 (
          nx2387), .B1 (nx2177)) ;
    inv01 ix2392 (.Y (nx2391), .A (A[12])) ;
    xnor2 ix1051 (.Y (nx1050), .A0 (nx2397), .A1 (nx1048)) ;
    nand02 ix2398 (.Y (nx2397), .A0 (nx3775), .A1 (nx3685)) ;
    xnor2 ix1049 (.Y (nx1048), .A0 (nx1032), .A1 (nx2403)) ;
    oai33 ix1033 (.Y (nx1032), .A0 (nx1627), .A1 (nx2165), .A2 (nx2185), .B0 (
          nx1631), .B1 (nx2391), .B2 (nx2189)) ;
    xnor2 ix2404 (.Y (nx2403), .A0 (nx2405), .A1 (nx2407)) ;
    nand02 ix2406 (.Y (nx2405), .A0 (nx3777), .A1 (nx3681)) ;
    xnor2 ix2408 (.Y (nx2407), .A0 (nx2409), .A1 (nx2411)) ;
    nand02 ix2410 (.Y (nx2409), .A0 (nx3781), .A1 (nx3677)) ;
    xnor2 ix2412 (.Y (nx2411), .A0 (nx2413), .A1 (nx2415)) ;
    nand02 ix2414 (.Y (nx2413), .A0 (nx3785), .A1 (nx3673)) ;
    nand02 ix2416 (.Y (nx2415), .A0 (nx3669), .A1 (nx3789)) ;
    nor02 ix939 (.Y (nx938), .A0 (nx2419), .A1 (nx2473)) ;
    nand02 ix2420 (.Y (nx2419), .A0 (nx662), .A1 (nx792)) ;
    nor02ii ix663 (.Y (nx662), .A0 (nx2423), .A1 (nx542)) ;
    xnor2 ix2424 (.Y (nx2423), .A0 (nx2205), .A1 (nx2289)) ;
    nor02 ix543 (.Y (nx542), .A0 (nx2427), .A1 (nx2469)) ;
    nand02 ix2428 (.Y (nx2427), .A0 (nx338), .A1 (nx432)) ;
    nor02ii ix339 (.Y (nx338), .A0 (nx2431), .A1 (nx254)) ;
    xnor2 ix2432 (.Y (nx2431), .A0 (nx2219), .A1 (nx2277)) ;
    nor02 ix255 (.Y (nx254), .A0 (nx2435), .A1 (nx2465)) ;
    nand02 ix2436 (.Y (nx2435), .A0 (nx122), .A1 (nx180)) ;
    nor02ii ix123 (.Y (nx122), .A0 (nx2439), .A1 (nx74)) ;
    xnor2 ix2440 (.Y (nx2439), .A0 (nx2233), .A1 (nx2265)) ;
    nor02 ix75 (.Y (nx74), .A0 (nx2443), .A1 (nx2461)) ;
    nand02 ix2444 (.Y (nx2443), .A0 (nx14), .A1 (nx36)) ;
    nor02 ix15 (.Y (nx14), .A0 (nx2447), .A1 (nx2451)) ;
    nand03 ix2448 (.Y (nx2447), .A0 (nx3785), .A1 (nx3723), .A2 (Product[0])) ;
    xnor2 ix2452 (.Y (nx2451), .A0 (nx2453), .A1 (nx2455)) ;
    nand02 ix2454 (.Y (nx2453), .A0 (nx3781), .A1 (nx3727)) ;
    xnor2 ix2456 (.Y (nx2455), .A0 (nx2253), .A1 (nx2255)) ;
    xnor2 ix37 (.Y (nx36), .A0 (nx20), .A1 (nx2257)) ;
    oai33 ix21 (.Y (nx20), .A0 (nx1627), .A1 (nx2195), .A2 (nx2455), .B0 (nx2253
          ), .B1 (nx1569), .B2 (nx1607)) ;
    xnor2 ix2462 (.Y (nx2461), .A0 (nx44), .A1 (nx70)) ;
    xnor2 ix181 (.Y (nx180), .A0 (nx128), .A1 (nx2269)) ;
    xnor2 ix2466 (.Y (nx2465), .A0 (nx188), .A1 (nx250)) ;
    xnor2 ix433 (.Y (nx432), .A0 (nx344), .A1 (nx2281)) ;
    xnor2 ix2470 (.Y (nx2469), .A0 (nx440), .A1 (nx538)) ;
    xnor2 ix793 (.Y (nx792), .A0 (nx668), .A1 (nx2293)) ;
    xnor2 ix2474 (.Y (nx2473), .A0 (nx800), .A1 (nx934)) ;
    xnor2 ix1261 (.Y (nx1260), .A0 (nx1100), .A1 (nx2481)) ;
    oai32 ix1101 (.Y (nx1100), .A0 (nx2479), .A1 (nx2195), .A2 (nx2305), .B0 (
          nx1553), .B1 (nx2301)) ;
    inv01 ix2480 (.Y (nx2479), .A (B[14])) ;
    xnor2 ix2482 (.Y (nx2481), .A0 (nx2483), .A1 (nx2485)) ;
    nand02 ix2484 (.Y (nx2483), .A0 (nx3729), .A1 (nx3727)) ;
    xnor2 ix2486 (.Y (nx2485), .A0 (nx2487), .A1 (nx2489)) ;
    aoi32 ix2488 (.Y (nx2487), .A0 (nx3737), .A1 (nx3723), .A2 (nx1084), .B0 (
          nx952), .B1 (nx1086)) ;
    xnor2 ix2490 (.Y (nx2489), .A0 (nx2491), .A1 (nx2493)) ;
    nand02 ix2492 (.Y (nx2491), .A0 (nx3733), .A1 (nx3723)) ;
    xnor2 ix2494 (.Y (nx2493), .A0 (nx1116), .A1 (nx1250)) ;
    oai32 ix1117 (.Y (nx1116), .A0 (nx2193), .A1 (nx1569), .A2 (nx2323), .B0 (
          nx2497), .B1 (nx2319)) ;
    inv01 ix2498 (.Y (nx2497), .A (nx960)) ;
    xnor2 ix1251 (.Y (nx1250), .A0 (nx2501), .A1 (nx1248)) ;
    nand02 ix2502 (.Y (nx2501), .A0 (nx3737), .A1 (nx3719)) ;
    xnor2 ix1249 (.Y (nx1248), .A0 (nx1124), .A1 (nx2507)) ;
    oai32 ix1125 (.Y (nx1124), .A0 (nx1559), .A1 (nx1733), .A2 (nx2331), .B0 (
          nx2325), .B1 (nx2327)) ;
    xnor2 ix2508 (.Y (nx2507), .A0 (nx2509), .A1 (nx2511)) ;
    nand02 ix2510 (.Y (nx2509), .A0 (nx3741), .A1 (nx3715)) ;
    xnor2 ix2512 (.Y (nx2511), .A0 (nx2513), .A1 (nx2515)) ;
    aoi32 ix2514 (.Y (nx2513), .A0 (nx3749), .A1 (nx3709), .A2 (nx1072), .B0 (
          nx976), .B1 (nx1074)) ;
    xnor2 ix2516 (.Y (nx2515), .A0 (nx2517), .A1 (nx2519)) ;
    nand02 ix2518 (.Y (nx2517), .A0 (nx3745), .A1 (nx3709)) ;
    xnor2 ix2520 (.Y (nx2519), .A0 (nx1140), .A1 (nx1238)) ;
    oai32 ix1141 (.Y (nx1140), .A0 (nx1567), .A1 (nx1589), .A2 (nx2349), .B0 (
          nx2523), .B1 (nx2345)) ;
    inv01 ix2524 (.Y (nx2523), .A (nx984)) ;
    xnor2 ix1239 (.Y (nx1238), .A0 (nx2527), .A1 (nx1236)) ;
    nand02 ix2528 (.Y (nx2527), .A0 (nx3749), .A1 (nx3705)) ;
    xnor2 ix1237 (.Y (nx1236), .A0 (nx1148), .A1 (nx2533)) ;
    oai32 ix1149 (.Y (nx1148), .A0 (nx1855), .A1 (nx1629), .A2 (nx2357), .B0 (
          nx2351), .B1 (nx2353)) ;
    xnor2 ix2534 (.Y (nx2533), .A0 (nx2535), .A1 (nx2537)) ;
    nand02 ix2536 (.Y (nx2535), .A0 (nx3753), .A1 (nx3701)) ;
    xnor2 ix2538 (.Y (nx2537), .A0 (nx2539), .A1 (nx2541)) ;
    aoi32 ix2540 (.Y (nx2539), .A0 (nx3763), .A1 (nx3697), .A2 (nx1060), .B0 (
          nx1000), .B1 (nx1062)) ;
    xnor2 ix2542 (.Y (nx2541), .A0 (nx2543), .A1 (nx2545)) ;
    nand02 ix2544 (.Y (nx2543), .A0 (nx3757), .A1 (nx3697)) ;
    xnor2 ix2546 (.Y (nx2545), .A0 (nx1164), .A1 (nx1226)) ;
    oai32 ix1165 (.Y (nx1164), .A0 (nx1731), .A1 (nx1703), .A2 (nx2375), .B0 (
          nx2549), .B1 (nx2371)) ;
    inv01 ix2550 (.Y (nx2549), .A (nx1008)) ;
    xnor2 ix1227 (.Y (nx1226), .A0 (nx2553), .A1 (nx1224)) ;
    nand02 ix2554 (.Y (nx2553), .A0 (nx3763), .A1 (nx3693)) ;
    xnor2 ix1225 (.Y (nx1224), .A0 (nx1172), .A1 (nx2559)) ;
    oai32 ix1173 (.Y (nx1172), .A0 (nx1579), .A1 (nx1825), .A2 (nx2383), .B0 (
          nx2377), .B1 (nx2379)) ;
    xnor2 ix2560 (.Y (nx2559), .A0 (nx2561), .A1 (nx2563)) ;
    nand02 ix2562 (.Y (nx2561), .A0 (nx3765), .A1 (nx3689)) ;
    xnor2 ix2564 (.Y (nx2563), .A0 (nx2565), .A1 (nx2567)) ;
    aoi32 ix2566 (.Y (nx2565), .A0 (nx3775), .A1 (nx3685), .A2 (nx1048), .B0 (
          nx1024), .B1 (nx1050)) ;
    xnor2 ix2568 (.Y (nx2567), .A0 (nx2569), .A1 (nx2571)) ;
    nand02 ix2570 (.Y (nx2569), .A0 (nx3769), .A1 (nx3685)) ;
    xnor2 ix2572 (.Y (nx2571), .A0 (nx1188), .A1 (nx1214)) ;
    oai32 ix1189 (.Y (nx1188), .A0 (nx1587), .A1 (nx2165), .A2 (nx2407), .B0 (
          nx2575), .B1 (nx2403)) ;
    inv01 ix2580 (.Y (nx2579), .A (A[13])) ;
    xnor2 ix1215 (.Y (nx1214), .A0 (nx2585), .A1 (nx1212)) ;
    nand02 ix2586 (.Y (nx2585), .A0 (nx3775), .A1 (nx3681)) ;
    xnor2 ix1213 (.Y (nx1212), .A0 (nx1196), .A1 (nx2591)) ;
    oai33 ix1197 (.Y (nx1196), .A0 (nx1627), .A1 (nx2391), .A2 (nx2411), .B0 (
          nx1631), .B1 (nx2579), .B2 (nx2415)) ;
    xnor2 ix2592 (.Y (nx2591), .A0 (nx2593), .A1 (nx2595)) ;
    nand02 ix2594 (.Y (nx2593), .A0 (nx3777), .A1 (nx3677)) ;
    xnor2 ix2596 (.Y (nx2595), .A0 (nx2597), .A1 (nx2599)) ;
    nand02 ix2598 (.Y (nx2597), .A0 (nx3781), .A1 (nx3673)) ;
    xnor2 ix2600 (.Y (nx2599), .A0 (nx2601), .A1 (nx2603)) ;
    nand02 ix2602 (.Y (nx2601), .A0 (nx3785), .A1 (nx3669)) ;
    nand02 ix2604 (.Y (nx2603), .A0 (nx3665), .A1 (nx3789)) ;
    nor02ii ix2879 (.Y (Product[1]), .A0 (nx2607), .A1 (nx2447)) ;
    aoi22 ix2608 (.Y (nx2607), .A0 (nx3723), .A1 (nx3789), .B0 (nx3787), .B1 (
          nx3727)) ;
    xor2 ix2869 (.Y (Product[2]), .A0 (nx2447), .A1 (nx2451)) ;
    xor2 ix2863 (.Y (Product[3]), .A0 (nx14), .A1 (nx36)) ;
    xor2 ix2857 (.Y (Product[4]), .A0 (nx2443), .A1 (nx2461)) ;
    xnor2 ix2851 (.Y (Product[5]), .A0 (nx74), .A1 (nx2439)) ;
    xor2 ix2845 (.Y (Product[6]), .A0 (nx122), .A1 (nx180)) ;
    xor2 ix2839 (.Y (Product[7]), .A0 (nx2435), .A1 (nx2465)) ;
    xnor2 ix2833 (.Y (Product[8]), .A0 (nx254), .A1 (nx2431)) ;
    xor2 ix2827 (.Y (Product[9]), .A0 (nx338), .A1 (nx432)) ;
    xor2 ix2821 (.Y (Product[10]), .A0 (nx2427), .A1 (nx2469)) ;
    xnor2 ix2815 (.Y (Product[11]), .A0 (nx542), .A1 (nx2423)) ;
    xor2 ix2809 (.Y (Product[12]), .A0 (nx662), .A1 (nx792)) ;
    xor2 ix2803 (.Y (Product[13]), .A0 (nx2419), .A1 (nx2473)) ;
    xnor2 ix2797 (.Y (Product[14]), .A0 (nx938), .A1 (nx1551)) ;
    xor2 ix2785 (.Y (Product[16]), .A0 (nx2637), .A1 (nx2639)) ;
    nand02 ix2638 (.Y (nx2637), .A0 (nx1094), .A1 (nx1260)) ;
    xnor2 ix2640 (.Y (nx2639), .A0 (nx1268), .A1 (nx1438)) ;
    oai32 ix1269 (.Y (nx1268), .A0 (nx2643), .A1 (nx2195), .A2 (nx2485), .B0 (
          nx2645), .B1 (nx2481)) ;
    inv01 ix2644 (.Y (nx2643), .A (B[15])) ;
    inv01 ix2646 (.Y (nx2645), .A (nx1100)) ;
    xnor2 ix1439 (.Y (nx1438), .A0 (nx1274), .A1 (nx2651)) ;
    oai32 ix1275 (.Y (nx1274), .A0 (nx2479), .A1 (nx1561), .A2 (nx2493), .B0 (
          nx2487), .B1 (nx2489)) ;
    xnor2 ix2652 (.Y (nx2651), .A0 (nx2653), .A1 (nx2655)) ;
    nand02 ix2654 (.Y (nx2653), .A0 (nx3729), .A1 (nx3723)) ;
    xnor2 ix2656 (.Y (nx2655), .A0 (nx2657), .A1 (nx2659)) ;
    aoi32 ix2658 (.Y (nx2657), .A0 (nx3737), .A1 (nx3719), .A2 (nx1248), .B0 (
          nx1116), .B1 (nx1250)) ;
    xnor2 ix2660 (.Y (nx2659), .A0 (nx2661), .A1 (nx2663)) ;
    nand02 ix2662 (.Y (nx2661), .A0 (nx3733), .A1 (nx3719)) ;
    xnor2 ix2664 (.Y (nx2663), .A0 (nx1290), .A1 (nx1428)) ;
    oai32 ix1291 (.Y (nx1290), .A0 (nx2193), .A1 (nx1733), .A2 (nx2511), .B0 (
          nx2667), .B1 (nx2507)) ;
    inv01 ix2668 (.Y (nx2667), .A (nx1124)) ;
    xnor2 ix1429 (.Y (nx1428), .A0 (nx2671), .A1 (nx1426)) ;
    nand02 ix2672 (.Y (nx2671), .A0 (nx3737), .A1 (nx3715)) ;
    xnor2 ix1427 (.Y (nx1426), .A0 (nx1298), .A1 (nx2677)) ;
    oai32 ix1299 (.Y (nx1298), .A0 (nx1559), .A1 (nx1581), .A2 (nx2519), .B0 (
          nx2513), .B1 (nx2515)) ;
    xnor2 ix2678 (.Y (nx2677), .A0 (nx2679), .A1 (nx2681)) ;
    nand02 ix2680 (.Y (nx2679), .A0 (nx3741), .A1 (nx3711)) ;
    xnor2 ix2682 (.Y (nx2681), .A0 (nx2683), .A1 (nx2685)) ;
    aoi32 ix2684 (.Y (nx2683), .A0 (nx3749), .A1 (nx3705), .A2 (nx1236), .B0 (
          nx1140), .B1 (nx1238)) ;
    xnor2 ix2686 (.Y (nx2685), .A0 (nx2687), .A1 (nx2689)) ;
    nand02 ix2688 (.Y (nx2687), .A0 (nx3745), .A1 (nx3705)) ;
    xnor2 ix2690 (.Y (nx2689), .A0 (nx1314), .A1 (nx1416)) ;
    oai32 ix1315 (.Y (nx1314), .A0 (nx1567), .A1 (nx1629), .A2 (nx2537), .B0 (
          nx2693), .B1 (nx2533)) ;
    inv01 ix2694 (.Y (nx2693), .A (nx1148)) ;
    xnor2 ix1417 (.Y (nx1416), .A0 (nx2697), .A1 (nx1414)) ;
    nand02 ix2698 (.Y (nx2697), .A0 (nx3749), .A1 (nx3701)) ;
    xnor2 ix1415 (.Y (nx1414), .A0 (nx1322), .A1 (nx2703)) ;
    oai32 ix1323 (.Y (nx1322), .A0 (nx1855), .A1 (nx1605), .A2 (nx2545), .B0 (
          nx2539), .B1 (nx2541)) ;
    xnor2 ix2704 (.Y (nx2703), .A0 (nx2705), .A1 (nx2707)) ;
    nand02 ix2706 (.Y (nx2705), .A0 (nx3753), .A1 (nx3697)) ;
    xnor2 ix2708 (.Y (nx2707), .A0 (nx2709), .A1 (nx2711)) ;
    aoi32 ix2710 (.Y (nx2709), .A0 (nx3763), .A1 (nx3693), .A2 (nx1224), .B0 (
          nx1164), .B1 (nx1226)) ;
    xnor2 ix2712 (.Y (nx2711), .A0 (nx2713), .A1 (nx2715)) ;
    nand02 ix2714 (.Y (nx2713), .A0 (nx3757), .A1 (nx3693)) ;
    xnor2 ix2716 (.Y (nx2715), .A0 (nx1338), .A1 (nx1404)) ;
    oai32 ix1339 (.Y (nx1338), .A0 (nx1731), .A1 (nx1825), .A2 (nx2563), .B0 (
          nx2719), .B1 (nx2559)) ;
    inv01 ix2720 (.Y (nx2719), .A (nx1172)) ;
    xnor2 ix1405 (.Y (nx1404), .A0 (nx2723), .A1 (nx1402)) ;
    nand02 ix2724 (.Y (nx2723), .A0 (nx3763), .A1 (nx3689)) ;
    xnor2 ix1403 (.Y (nx1402), .A0 (nx1346), .A1 (nx2729)) ;
    oai32 ix1347 (.Y (nx1346), .A0 (nx1579), .A1 (nx1979), .A2 (nx2571), .B0 (
          nx2565), .B1 (nx2567)) ;
    xnor2 ix2730 (.Y (nx2729), .A0 (nx2731), .A1 (nx2733)) ;
    nand02 ix2732 (.Y (nx2731), .A0 (nx3765), .A1 (nx3685)) ;
    xnor2 ix2734 (.Y (nx2733), .A0 (nx2735), .A1 (nx2737)) ;
    aoi32 ix2736 (.Y (nx2735), .A0 (nx3775), .A1 (nx3681), .A2 (nx1212), .B0 (
          nx1188), .B1 (nx1214)) ;
    xnor2 ix2738 (.Y (nx2737), .A0 (nx2739), .A1 (nx2741)) ;
    nand02 ix2740 (.Y (nx2739), .A0 (nx3769), .A1 (nx3681)) ;
    xnor2 ix2742 (.Y (nx2741), .A0 (nx1362), .A1 (nx1392)) ;
    oai32 ix1363 (.Y (nx1362), .A0 (nx1587), .A1 (nx2391), .A2 (nx2595), .B0 (
          nx2745), .B1 (nx2591)) ;
    inv01 ix2750 (.Y (nx2749), .A (A[14])) ;
    xnor2 ix1393 (.Y (nx1392), .A0 (nx2755), .A1 (nx1390)) ;
    nand02 ix2756 (.Y (nx2755), .A0 (nx3775), .A1 (nx3677)) ;
    xnor2 ix1391 (.Y (nx1390), .A0 (nx1370), .A1 (nx2763)) ;
    oai33 ix1371 (.Y (nx1370), .A0 (nx1627), .A1 (nx2579), .A2 (nx2599), .B0 (
          nx2601), .B1 (nx2761), .B2 (nx1607)) ;
    inv01 ix2762 (.Y (nx2761), .A (A[15])) ;
    xnor2 ix2764 (.Y (nx2763), .A0 (nx2765), .A1 (nx2767)) ;
    nand02 ix2766 (.Y (nx2765), .A0 (nx3777), .A1 (nx3673)) ;
    nand02 ix2768 (.Y (nx2767), .A0 (nx2769), .A1 (nx1382)) ;
    nand04 ix2770 (.Y (nx2769), .A0 (nx3781), .A1 (nx3665), .A2 (nx3787), .A3 (
           nx3669)) ;
    xnor2 ix2783 (.Y (Product[17]), .A0 (nx2775), .A1 (nx1604)) ;
    aoi22 ix2776 (.Y (nx2775), .A0 (nx1268), .A1 (nx1438), .B0 (nx1262), .B1 (
          nx1440)) ;
    xnor2 ix1605 (.Y (nx1604), .A0 (nx1452), .A1 (nx2787)) ;
    oai32 ix1453 (.Y (nx1452), .A0 (nx2643), .A1 (nx1561), .A2 (nx2655), .B0 (
          nx2785), .B1 (nx2651)) ;
    inv01 ix2786 (.Y (nx2785), .A (nx1274)) ;
    xnor2 ix2788 (.Y (nx2787), .A0 (nx1458), .A1 (nx1600)) ;
    oai32 ix1459 (.Y (nx1458), .A0 (nx2479), .A1 (nx1569), .A2 (nx2663), .B0 (
          nx2657), .B1 (nx2659)) ;
    xnor2 ix1601 (.Y (nx1600), .A0 (nx2793), .A1 (nx1598)) ;
    nand02 ix2794 (.Y (nx2793), .A0 (nx3729), .A1 (nx3719)) ;
    xnor2 ix1599 (.Y (nx1598), .A0 (nx2797), .A1 (nx1596)) ;
    aoi32 ix2798 (.Y (nx2797), .A0 (nx3737), .A1 (nx3715), .A2 (nx1426), .B0 (
          nx1290), .B1 (nx1428)) ;
    xnor2 ix1597 (.Y (nx1596), .A0 (nx2801), .A1 (nx1594)) ;
    nand02 ix2802 (.Y (nx2801), .A0 (nx3733), .A1 (nx3715)) ;
    xnor2 ix1595 (.Y (nx1594), .A0 (nx1474), .A1 (nx2809)) ;
    oai32 ix1475 (.Y (nx1474), .A0 (nx2193), .A1 (nx1581), .A2 (nx2681), .B0 (
          nx2807), .B1 (nx2677)) ;
    inv01 ix2808 (.Y (nx2807), .A (nx1298)) ;
    xnor2 ix2810 (.Y (nx2809), .A0 (nx2811), .A1 (nx2813)) ;
    nand02 ix2812 (.Y (nx2811), .A0 (nx3737), .A1 (nx3711)) ;
    xnor2 ix2814 (.Y (nx2813), .A0 (nx1482), .A1 (nx1588)) ;
    oai32 ix1483 (.Y (nx1482), .A0 (nx1559), .A1 (nx1589), .A2 (nx2689), .B0 (
          nx2683), .B1 (nx2685)) ;
    xnor2 ix1589 (.Y (nx1588), .A0 (nx2819), .A1 (nx1586)) ;
    nand02 ix2820 (.Y (nx2819), .A0 (nx3741), .A1 (nx3707)) ;
    xnor2 ix1587 (.Y (nx1586), .A0 (nx2823), .A1 (nx1584)) ;
    aoi32 ix2824 (.Y (nx2823), .A0 (nx3749), .A1 (nx3701), .A2 (nx1414), .B0 (
          nx1314), .B1 (nx1416)) ;
    xnor2 ix1585 (.Y (nx1584), .A0 (nx2827), .A1 (nx1582)) ;
    nand02 ix2828 (.Y (nx2827), .A0 (nx3745), .A1 (nx3701)) ;
    xnor2 ix1583 (.Y (nx1582), .A0 (nx1498), .A1 (nx2835)) ;
    oai32 ix1499 (.Y (nx1498), .A0 (nx1567), .A1 (nx1605), .A2 (nx2707), .B0 (
          nx2833), .B1 (nx2703)) ;
    inv01 ix2834 (.Y (nx2833), .A (nx1322)) ;
    xnor2 ix2836 (.Y (nx2835), .A0 (nx2837), .A1 (nx2839)) ;
    nand02 ix2838 (.Y (nx2837), .A0 (nx3749), .A1 (nx3697)) ;
    xnor2 ix2840 (.Y (nx2839), .A0 (nx1506), .A1 (nx1576)) ;
    oai32 ix1507 (.Y (nx1506), .A0 (nx1855), .A1 (nx1703), .A2 (nx2715), .B0 (
          nx2709), .B1 (nx2711)) ;
    xnor2 ix1577 (.Y (nx1576), .A0 (nx2845), .A1 (nx1574)) ;
    nand02 ix2846 (.Y (nx2845), .A0 (nx3753), .A1 (nx3693)) ;
    xnor2 ix1575 (.Y (nx1574), .A0 (nx2849), .A1 (nx1572)) ;
    aoi32 ix2850 (.Y (nx2849), .A0 (nx3763), .A1 (nx3689), .A2 (nx1402), .B0 (
          nx1338), .B1 (nx1404)) ;
    xnor2 ix1573 (.Y (nx1572), .A0 (nx2853), .A1 (nx1570)) ;
    nand02 ix2854 (.Y (nx2853), .A0 (nx3757), .A1 (nx3689)) ;
    xnor2 ix1571 (.Y (nx1570), .A0 (nx1522), .A1 (nx2861)) ;
    oai32 ix1523 (.Y (nx1522), .A0 (nx1731), .A1 (nx1979), .A2 (nx2733), .B0 (
          nx2859), .B1 (nx2729)) ;
    inv01 ix2860 (.Y (nx2859), .A (nx1346)) ;
    xnor2 ix2862 (.Y (nx2861), .A0 (nx2863), .A1 (nx2865)) ;
    nand02 ix2864 (.Y (nx2863), .A0 (nx3763), .A1 (nx3685)) ;
    xnor2 ix2866 (.Y (nx2865), .A0 (nx1530), .A1 (nx1564)) ;
    oai32 ix1531 (.Y (nx1530), .A0 (nx1579), .A1 (nx2165), .A2 (nx2741), .B0 (
          nx2735), .B1 (nx2737)) ;
    xnor2 ix1565 (.Y (nx1564), .A0 (nx2871), .A1 (nx1562)) ;
    nand02 ix2872 (.Y (nx2871), .A0 (nx3765), .A1 (nx3681)) ;
    xnor2 ix1563 (.Y (nx1562), .A0 (nx2875), .A1 (nx1560)) ;
    aoi32 ix2876 (.Y (nx2875), .A0 (nx3775), .A1 (nx3677), .A2 (nx1390), .B0 (
          nx1362), .B1 (nx1392)) ;
    xnor2 ix1561 (.Y (nx1560), .A0 (nx2879), .A1 (nx1558)) ;
    nand02 ix2880 (.Y (nx2879), .A0 (nx3769), .A1 (nx3677)) ;
    xnor2 ix1559 (.Y (nx1558), .A0 (nx1546), .A1 (nx2887)) ;
    oai32 ix1547 (.Y (nx1546), .A0 (nx1587), .A1 (nx2579), .A2 (nx2767), .B0 (
          nx2883), .B1 (nx2763)) ;
    xnor2 ix2888 (.Y (nx2887), .A0 (nx2889), .A1 (nx2891)) ;
    nand02 ix2890 (.Y (nx2889), .A0 (nx3775), .A1 (nx3673)) ;
    xnor2 ix2892 (.Y (nx2891), .A0 (nx2769), .A1 (nx2893)) ;
    xnor2 ix2894 (.Y (nx2893), .A0 (nx2895), .A1 (nx2897)) ;
    nand02 ix2896 (.Y (nx2895), .A0 (nx3777), .A1 (nx3669)) ;
    nand02 ix2898 (.Y (nx2897), .A0 (nx3783), .A1 (nx3665)) ;
    xnor2 ix2781 (.Y (Product[18]), .A0 (nx2900), .A1 (nx1764)) ;
    aoi22 ix2901 (.Y (nx2900), .A0 (nx1452), .A1 (nx1602), .B0 (nx1446), .B1 (
          nx1604)) ;
    xnor2 ix1765 (.Y (nx1764), .A0 (nx2907), .A1 (nx1762)) ;
    aoi32 ix2908 (.Y (nx2907), .A0 (nx3729), .A1 (nx3719), .A2 (nx1598), .B0 (
          nx1458), .B1 (nx1600)) ;
    xnor2 ix1763 (.Y (nx1762), .A0 (nx2910), .A1 (nx1760)) ;
    aoi32 ix2911 (.Y (nx2910), .A0 (nx3733), .A1 (nx3715), .A2 (nx1594), .B0 (
          nx1466), .B1 (nx1596)) ;
    xnor2 ix1761 (.Y (nx1760), .A0 (nx2914), .A1 (nx1758)) ;
    nand02 ix2915 (.Y (nx2914), .A0 (nx3729), .A1 (nx3715)) ;
    xnor2 ix1759 (.Y (nx1758), .A0 (nx1630), .A1 (nx2924)) ;
    oai32 ix1631 (.Y (nx1630), .A0 (nx2918), .A1 (nx1581), .A2 (nx2813), .B0 (
          nx2920), .B1 (nx2809)) ;
    inv01 ix2919 (.Y (nx2918), .A (B[13])) ;
    xnor2 ix2925 (.Y (nx2924), .A0 (nx2926), .A1 (nx2928)) ;
    nand02 ix2927 (.Y (nx2926), .A0 (nx3733), .A1 (nx3711)) ;
    xnor2 ix2929 (.Y (nx2928), .A0 (nx2930), .A1 (nx2932)) ;
    aoi32 ix2931 (.Y (nx2930), .A0 (nx3741), .A1 (nx3707), .A2 (nx1586), .B0 (
          nx1482), .B1 (nx1588)) ;
    xnor2 ix2933 (.Y (nx2932), .A0 (nx2934), .A1 (nx2936)) ;
    nand02 ix2935 (.Y (nx2934), .A0 (nx3737), .A1 (nx3707)) ;
    xnor2 ix2937 (.Y (nx2936), .A0 (nx2938), .A1 (nx2941)) ;
    aoi32 ix2939 (.Y (nx2938), .A0 (nx3745), .A1 (nx3703), .A2 (nx1582), .B0 (
          nx1490), .B1 (nx1584)) ;
    xnor2 ix2942 (.Y (nx2941), .A0 (nx2943), .A1 (nx2945)) ;
    nand02 ix2944 (.Y (nx2943), .A0 (nx3741), .A1 (nx3703)) ;
    xnor2 ix2946 (.Y (nx2945), .A0 (nx1654), .A1 (nx1744)) ;
    oai32 ix1655 (.Y (nx1654), .A0 (nx2948), .A1 (nx1605), .A2 (nx2839), .B0 (
          nx2950), .B1 (nx2835)) ;
    inv01 ix2949 (.Y (nx2948), .A (B[10])) ;
    xnor2 ix1745 (.Y (nx1744), .A0 (nx2955), .A1 (nx1742)) ;
    nand02 ix2956 (.Y (nx2955), .A0 (nx3745), .A1 (nx3697)) ;
    xnor2 ix1743 (.Y (nx1742), .A0 (nx2958), .A1 (nx1740)) ;
    aoi32 ix2959 (.Y (nx2958), .A0 (nx3753), .A1 (nx3693), .A2 (nx1574), .B0 (
          nx1506), .B1 (nx1576)) ;
    xnor2 ix1741 (.Y (nx1740), .A0 (nx2961), .A1 (nx1738)) ;
    nand02 ix2962 (.Y (nx2961), .A0 (nx3751), .A1 (nx3693)) ;
    xnor2 ix1739 (.Y (nx1738), .A0 (nx2964), .A1 (nx1736)) ;
    aoi32 ix2965 (.Y (nx2964), .A0 (nx3757), .A1 (nx3689), .A2 (nx1570), .B0 (
          nx1514), .B1 (nx1572)) ;
    xnor2 ix1737 (.Y (nx1736), .A0 (nx2968), .A1 (nx1734)) ;
    nand02 ix2969 (.Y (nx2968), .A0 (nx3753), .A1 (nx3689)) ;
    xnor2 ix1735 (.Y (nx1734), .A0 (nx1678), .A1 (nx2978)) ;
    oai32 ix1679 (.Y (nx1678), .A0 (nx2972), .A1 (nx1979), .A2 (nx2865), .B0 (
          nx2974), .B1 (nx2861)) ;
    inv01 ix2973 (.Y (nx2972), .A (B[7])) ;
    xnor2 ix2979 (.Y (nx2978), .A0 (nx2980), .A1 (nx2982)) ;
    nand02 ix2981 (.Y (nx2980), .A0 (nx3757), .A1 (nx3685)) ;
    xnor2 ix2983 (.Y (nx2982), .A0 (nx2984), .A1 (nx2986)) ;
    aoi32 ix2985 (.Y (nx2984), .A0 (nx3765), .A1 (nx3681), .A2 (nx1562), .B0 (
          nx1530), .B1 (nx1564)) ;
    xnor2 ix2987 (.Y (nx2986), .A0 (nx2988), .A1 (nx2990)) ;
    nand02 ix2989 (.Y (nx2988), .A0 (nx3763), .A1 (nx3681)) ;
    xnor2 ix2991 (.Y (nx2990), .A0 (nx2992), .A1 (nx2995)) ;
    aoi32 ix2993 (.Y (nx2992), .A0 (nx3769), .A1 (nx3677), .A2 (nx1558), .B0 (
          nx1538), .B1 (nx1560)) ;
    xnor2 ix2996 (.Y (nx2995), .A0 (nx2997), .A1 (nx2999)) ;
    nand02 ix2998 (.Y (nx2997), .A0 (nx3765), .A1 (nx3677)) ;
    xnor2 ix3000 (.Y (nx2999), .A0 (nx1702), .A1 (nx1720)) ;
    oai32 ix1703 (.Y (nx1702), .A0 (nx3002), .A1 (nx2579), .A2 (nx2891), .B0 (
          nx3004), .B1 (nx2887)) ;
    inv01 ix3003 (.Y (nx3002), .A (B[4])) ;
    aoi22 ix3008 (.Y (nx3007), .A0 (nx3787), .A1 (nx3665), .B0 (nx3783), .B1 (
          nx3669)) ;
    xnor2 ix1721 (.Y (nx1720), .A0 (nx3011), .A1 (nx1718)) ;
    nand02 ix3012 (.Y (nx3011), .A0 (nx3769), .A1 (nx3673)) ;
    xnor2 ix1719 (.Y (nx1718), .A0 (nx1710), .A1 (nx3015)) ;
    aoi21 ix1711 (.Y (nx1710), .A0 (nx2895), .A1 (nx2601), .B0 (nx2897)) ;
    xnor2 ix3016 (.Y (nx3015), .A0 (nx3017), .A1 (nx3019)) ;
    nand02 ix3018 (.Y (nx3017), .A0 (nx3775), .A1 (nx3669)) ;
    nand02 ix3020 (.Y (nx3019), .A0 (nx3779), .A1 (nx3665)) ;
    xor2 ix2779 (.Y (Product[19]), .A0 (nx1770), .A1 (nx1912)) ;
    oai22 ix1771 (.Y (nx1770), .A0 (nx2900), .A1 (nx3023), .B0 (nx2907), .B1 (
          nx3025)) ;
    xnor2 ix1913 (.Y (nx1912), .A0 (nx3028), .A1 (nx1910)) ;
    aoi32 ix3029 (.Y (nx3028), .A0 (nx3729), .A1 (nx3715), .A2 (nx1758), .B0 (
          nx1622), .B1 (nx1760)) ;
    xnor2 ix1911 (.Y (nx1910), .A0 (nx1782), .A1 (nx3037)) ;
    oai32 ix1783 (.Y (nx1782), .A0 (nx2479), .A1 (nx1581), .A2 (nx2928), .B0 (
          nx3033), .B1 (nx2924)) ;
    xnor2 ix3038 (.Y (nx3037), .A0 (nx3039), .A1 (nx3041)) ;
    nand02 ix3040 (.Y (nx3039), .A0 (nx3729), .A1 (nx3711)) ;
    xnor2 ix3042 (.Y (nx3041), .A0 (nx1790), .A1 (nx1904)) ;
    oai32 ix1791 (.Y (nx1790), .A0 (nx2918), .A1 (nx1589), .A2 (nx2936), .B0 (
          nx2930), .B1 (nx2932)) ;
    xnor2 ix1905 (.Y (nx1904), .A0 (nx3045), .A1 (nx1902)) ;
    nand02 ix3046 (.Y (nx3045), .A0 (nx3733), .A1 (nx3707)) ;
    xnor2 ix1903 (.Y (nx1902), .A0 (nx1798), .A1 (nx3049)) ;
    oai32 ix1799 (.Y (nx1798), .A0 (nx2193), .A1 (nx1629), .A2 (nx2945), .B0 (
          nx2938), .B1 (nx2941)) ;
    xnor2 ix3050 (.Y (nx3049), .A0 (nx3051), .A1 (nx3053)) ;
    nand02 ix3052 (.Y (nx3051), .A0 (nx3737), .A1 (nx3703)) ;
    xnor2 ix3054 (.Y (nx3053), .A0 (nx3055), .A1 (nx3057)) ;
    aoi32 ix3056 (.Y (nx3055), .A0 (nx3745), .A1 (nx3697), .A2 (nx1742), .B0 (
          nx1654), .B1 (nx1744)) ;
    xnor2 ix3058 (.Y (nx3057), .A0 (nx3059), .A1 (nx3061)) ;
    nand02 ix3060 (.Y (nx3059), .A0 (nx3741), .A1 (nx3699)) ;
    xnor2 ix3062 (.Y (nx3061), .A0 (nx3063), .A1 (nx3066)) ;
    aoi32 ix3064 (.Y (nx3063), .A0 (nx3751), .A1 (nx3693), .A2 (nx1738), .B0 (
          nx1662), .B1 (nx1740)) ;
    xnor2 ix3067 (.Y (nx3066), .A0 (nx3068), .A1 (nx3070)) ;
    nand02 ix3069 (.Y (nx3068), .A0 (nx3745), .A1 (nx3695)) ;
    xnor2 ix3071 (.Y (nx3070), .A0 (nx3072), .A1 (nx3075)) ;
    aoi32 ix3073 (.Y (nx3072), .A0 (nx3753), .A1 (nx3689), .A2 (nx1734), .B0 (
          nx1670), .B1 (nx1736)) ;
    xnor2 ix3076 (.Y (nx3075), .A0 (nx3077), .A1 (nx3079)) ;
    nand02 ix3078 (.Y (nx3077), .A0 (nx3751), .A1 (nx3689)) ;
    xnor2 ix3080 (.Y (nx3079), .A0 (nx1830), .A1 (nx1884)) ;
    oai32 ix1831 (.Y (nx1830), .A0 (nx1855), .A1 (nx1979), .A2 (nx2982), .B0 (
          nx3082), .B1 (nx2978)) ;
    xnor2 ix1885 (.Y (nx1884), .A0 (nx3087), .A1 (nx1882)) ;
    nand02 ix3088 (.Y (nx3087), .A0 (nx3753), .A1 (nx3685)) ;
    xnor2 ix1883 (.Y (nx1882), .A0 (nx1838), .A1 (nx3091)) ;
    oai32 ix1839 (.Y (nx1838), .A0 (nx2972), .A1 (nx2165), .A2 (nx2990), .B0 (
          nx2984), .B1 (nx2986)) ;
    xnor2 ix3092 (.Y (nx3091), .A0 (nx3093), .A1 (nx3095)) ;
    nand02 ix3094 (.Y (nx3093), .A0 (nx3757), .A1 (nx3681)) ;
    xnor2 ix3096 (.Y (nx3095), .A0 (nx1846), .A1 (nx1876)) ;
    oai32 ix1847 (.Y (nx1846), .A0 (nx1731), .A1 (nx2391), .A2 (nx2999), .B0 (
          nx2992), .B1 (nx2995)) ;
    xnor2 ix1877 (.Y (nx1876), .A0 (nx3099), .A1 (nx1874)) ;
    nand02 ix3100 (.Y (nx3099), .A0 (nx3763), .A1 (nx3677)) ;
    xnor2 ix1875 (.Y (nx1874), .A0 (nx3102), .A1 (nx1872)) ;
    aoi32 ix3103 (.Y (nx3102), .A0 (nx3771), .A1 (nx3673), .A2 (nx1718), .B0 (
          nx1702), .B1 (nx1720)) ;
    xnor2 ix1873 (.Y (nx1872), .A0 (nx3105), .A1 (nx1870)) ;
    nand02 ix3106 (.Y (nx3105), .A0 (nx3765), .A1 (nx3673)) ;
    xnor2 ix1871 (.Y (nx1870), .A0 (nx1862), .A1 (nx3111)) ;
    oai32 ix1863 (.Y (nx1862), .A0 (nx3002), .A1 (nx2749), .A2 (nx3019), .B0 (
          nx3109), .B1 (nx3015)) ;
    xnor2 ix3112 (.Y (nx3111), .A0 (nx3113), .A1 (nx3115)) ;
    nand02 ix3114 (.Y (nx3113), .A0 (nx3771), .A1 (nx3669)) ;
    nand02 ix3116 (.Y (nx3115), .A0 (nx3775), .A1 (nx3665)) ;
    xnor2 ix2777 (.Y (Product[20]), .A0 (nx3118), .A1 (nx2048)) ;
    aoi22 ix3119 (.Y (nx3118), .A0 (nx1776), .A1 (nx1910), .B0 (nx1770), .B1 (
          nx1912)) ;
    xnor2 ix2049 (.Y (nx2048), .A0 (nx1924), .A1 (nx3127)) ;
    oai32 ix1925 (.Y (nx1924), .A0 (nx2643), .A1 (nx1581), .A2 (nx3041), .B0 (
          nx3123), .B1 (nx3037)) ;
    xnor2 ix3128 (.Y (nx3127), .A0 (nx3129), .A1 (nx3131)) ;
    aoi32 ix3130 (.Y (nx3129), .A0 (nx3733), .A1 (nx3707), .A2 (nx1902), .B0 (
          nx1790), .B1 (nx1904)) ;
    xnor2 ix3132 (.Y (nx3131), .A0 (nx3133), .A1 (nx3135)) ;
    nand02 ix3134 (.Y (nx3133), .A0 (nx3729), .A1 (nx3707)) ;
    xnor2 ix3136 (.Y (nx3135), .A0 (nx1938), .A1 (nx2040)) ;
    oai32 ix1939 (.Y (nx1938), .A0 (nx2918), .A1 (nx1629), .A2 (nx3053), .B0 (
          nx3138), .B1 (nx3049)) ;
    inv01 ix3139 (.Y (nx3138), .A (nx1798)) ;
    xnor2 ix2041 (.Y (nx2040), .A0 (nx3141), .A1 (nx2038)) ;
    nand02 ix3142 (.Y (nx3141), .A0 (nx3733), .A1 (nx3703)) ;
    xnor2 ix2039 (.Y (nx2038), .A0 (nx1946), .A1 (nx3145)) ;
    oai32 ix1947 (.Y (nx1946), .A0 (nx2193), .A1 (nx1605), .A2 (nx3061), .B0 (
          nx3055), .B1 (nx3057)) ;
    xnor2 ix3146 (.Y (nx3145), .A0 (nx3147), .A1 (nx3149)) ;
    nand02 ix3148 (.Y (nx3147), .A0 (nx3737), .A1 (nx3699)) ;
    xnor2 ix3150 (.Y (nx3149), .A0 (nx1954), .A1 (nx2032)) ;
    oai32 ix1955 (.Y (nx1954), .A0 (nx1559), .A1 (nx1703), .A2 (nx3070), .B0 (
          nx3063), .B1 (nx3066)) ;
    xnor2 ix2033 (.Y (nx2032), .A0 (nx3153), .A1 (nx2030)) ;
    nand02 ix3154 (.Y (nx3153), .A0 (nx3741), .A1 (nx3695)) ;
    xnor2 ix2031 (.Y (nx2030), .A0 (nx1962), .A1 (nx3157)) ;
    oai32 ix1963 (.Y (nx1962), .A0 (nx2948), .A1 (nx1825), .A2 (nx3079), .B0 (
          nx3072), .B1 (nx3075)) ;
    xnor2 ix3158 (.Y (nx3157), .A0 (nx3159), .A1 (nx3161)) ;
    nand02 ix3160 (.Y (nx3159), .A0 (nx3745), .A1 (nx3691)) ;
    xnor2 ix3162 (.Y (nx3161), .A0 (nx3163), .A1 (nx3165)) ;
    aoi32 ix3164 (.Y (nx3163), .A0 (nx3753), .A1 (nx3685), .A2 (nx1882), .B0 (
          nx1830), .B1 (nx1884)) ;
    xnor2 ix3166 (.Y (nx3165), .A0 (nx3167), .A1 (nx3169)) ;
    nand02 ix3168 (.Y (nx3167), .A0 (nx3751), .A1 (nx3685)) ;
    xnor2 ix3170 (.Y (nx3169), .A0 (nx1978), .A1 (nx2020)) ;
    oai32 ix1979 (.Y (nx1978), .A0 (nx1855), .A1 (nx2165), .A2 (nx3095), .B0 (
          nx3172), .B1 (nx3091)) ;
    inv01 ix3173 (.Y (nx3172), .A (nx1838)) ;
    xnor2 ix2021 (.Y (nx2020), .A0 (nx3175), .A1 (nx2018)) ;
    nand02 ix3176 (.Y (nx3175), .A0 (nx3753), .A1 (nx3681)) ;
    xnor2 ix2019 (.Y (nx2018), .A0 (nx3178), .A1 (nx2016)) ;
    aoi32 ix3179 (.Y (nx3178), .A0 (nx3763), .A1 (nx3677), .A2 (nx1874), .B0 (
          nx1846), .B1 (nx1876)) ;
    xnor2 ix2017 (.Y (nx2016), .A0 (nx3181), .A1 (nx2014)) ;
    nand02 ix3182 (.Y (nx3181), .A0 (nx3757), .A1 (nx3677)) ;
    xnor2 ix2015 (.Y (nx2014), .A0 (nx3184), .A1 (nx2012)) ;
    aoi32 ix3185 (.Y (nx3184), .A0 (nx3767), .A1 (nx3673), .A2 (nx1870), .B0 (
          nx1854), .B1 (nx1872)) ;
    xnor2 ix2013 (.Y (nx2012), .A0 (nx3188), .A1 (nx2010)) ;
    nand02 ix3189 (.Y (nx3188), .A0 (nx3763), .A1 (nx3673)) ;
    xnor2 ix2011 (.Y (nx2010), .A0 (nx2002), .A1 (nx3196)) ;
    oai32 ix2003 (.Y (nx2002), .A0 (nx1579), .A1 (nx2749), .A2 (nx3115), .B0 (
          nx3192), .B1 (nx3111)) ;
    xnor2 ix3197 (.Y (nx3196), .A0 (nx3198), .A1 (nx3200)) ;
    nand02 ix3199 (.Y (nx3198), .A0 (nx3767), .A1 (nx3669)) ;
    nand02 ix3201 (.Y (nx3200), .A0 (nx3771), .A1 (nx3665)) ;
    xor2 ix2775 (.Y (Product[21]), .A0 (nx2054), .A1 (nx2172)) ;
    oai22 ix2055 (.Y (nx2054), .A0 (nx3118), .A1 (nx3204), .B0 (nx3206), .B1 (
          nx3127)) ;
    xnor2 ix2173 (.Y (nx2172), .A0 (nx2060), .A1 (nx3212)) ;
    oai32 ix2061 (.Y (nx2060), .A0 (nx2643), .A1 (nx1589), .A2 (nx3135), .B0 (
          nx3129), .B1 (nx3131)) ;
    xnor2 ix3213 (.Y (nx3212), .A0 (nx3214), .A1 (nx3216)) ;
    aoi32 ix3215 (.Y (nx3214), .A0 (nx3733), .A1 (nx3703), .A2 (nx2038), .B0 (
          nx1938), .B1 (nx2040)) ;
    xnor2 ix3217 (.Y (nx3216), .A0 (nx3218), .A1 (nx3220)) ;
    nand02 ix3219 (.Y (nx3218), .A0 (nx3729), .A1 (nx3703)) ;
    xnor2 ix3221 (.Y (nx3220), .A0 (nx2074), .A1 (nx2164)) ;
    oai32 ix2075 (.Y (nx2074), .A0 (nx2918), .A1 (nx1605), .A2 (nx3149), .B0 (
          nx3223), .B1 (nx3145)) ;
    inv01 ix3224 (.Y (nx3223), .A (nx1946)) ;
    xnor2 ix2165 (.Y (nx2164), .A0 (nx3226), .A1 (nx2162)) ;
    nand02 ix3227 (.Y (nx3226), .A0 (nx3733), .A1 (nx3699)) ;
    xnor2 ix2163 (.Y (nx2162), .A0 (nx3229), .A1 (nx2160)) ;
    aoi32 ix3230 (.Y (nx3229), .A0 (nx3741), .A1 (nx3695), .A2 (nx2030), .B0 (
          nx1954), .B1 (nx2032)) ;
    xnor2 ix2161 (.Y (nx2160), .A0 (nx3232), .A1 (nx2158)) ;
    nand02 ix3233 (.Y (nx3232), .A0 (nx3737), .A1 (nx3695)) ;
    xnor2 ix2159 (.Y (nx2158), .A0 (nx2090), .A1 (nx3238)) ;
    oai32 ix2091 (.Y (nx2090), .A0 (nx1559), .A1 (nx1825), .A2 (nx3161), .B0 (
          nx3236), .B1 (nx3157)) ;
    inv01 ix3237 (.Y (nx3236), .A (nx1962)) ;
    xnor2 ix3239 (.Y (nx3238), .A0 (nx3240), .A1 (nx3242)) ;
    nand02 ix3241 (.Y (nx3240), .A0 (nx3741), .A1 (nx3691)) ;
    xnor2 ix3243 (.Y (nx3242), .A0 (nx2098), .A1 (nx2152)) ;
    oai32 ix2099 (.Y (nx2098), .A0 (nx2948), .A1 (nx1979), .A2 (nx3169), .B0 (
          nx3163), .B1 (nx3165)) ;
    xnor2 ix2153 (.Y (nx2152), .A0 (nx3246), .A1 (nx2150)) ;
    nand02 ix3247 (.Y (nx3246), .A0 (nx3745), .A1 (nx3685)) ;
    xnor2 ix2151 (.Y (nx2150), .A0 (nx3249), .A1 (nx2148)) ;
    aoi32 ix3250 (.Y (nx3249), .A0 (nx3755), .A1 (nx3681), .A2 (nx2018), .B0 (
          nx1978), .B1 (nx2020)) ;
    xnor2 ix2149 (.Y (nx2148), .A0 (nx3252), .A1 (nx2146)) ;
    nand02 ix3253 (.Y (nx3252), .A0 (nx3751), .A1 (nx3681)) ;
    xnor2 ix2147 (.Y (nx2146), .A0 (nx3255), .A1 (nx2144)) ;
    aoi32 ix3256 (.Y (nx3255), .A0 (nx3757), .A1 (nx3677), .A2 (nx2014), .B0 (
          nx1986), .B1 (nx2016)) ;
    xnor2 ix2145 (.Y (nx2144), .A0 (nx3259), .A1 (nx2142)) ;
    nand02 ix3260 (.Y (nx3259), .A0 (nx3755), .A1 (nx3677)) ;
    xnor2 ix2143 (.Y (nx2142), .A0 (nx3262), .A1 (nx2140)) ;
    aoi32 ix3263 (.Y (nx3262), .A0 (nx3763), .A1 (nx3673), .A2 (nx2010), .B0 (
          nx1994), .B1 (nx2012)) ;
    xnor2 ix2141 (.Y (nx2140), .A0 (nx3266), .A1 (nx2138)) ;
    nand02 ix3267 (.Y (nx3266), .A0 (nx3759), .A1 (nx3673)) ;
    xnor2 ix2139 (.Y (nx2138), .A0 (nx2130), .A1 (nx3274)) ;
    oai32 ix2131 (.Y (nx2130), .A0 (nx1731), .A1 (nx2749), .A2 (nx3200), .B0 (
          nx3270), .B1 (nx3196)) ;
    xnor2 ix3275 (.Y (nx3274), .A0 (nx3276), .A1 (nx3278)) ;
    nand02 ix3277 (.Y (nx3276), .A0 (nx3763), .A1 (nx3669)) ;
    nand02 ix3279 (.Y (nx3278), .A0 (nx3767), .A1 (nx3665)) ;
    xnor2 ix2773 (.Y (Product[22]), .A0 (nx3281), .A1 (nx2284)) ;
    aoi22 ix3282 (.Y (nx3281), .A0 (nx2060), .A1 (nx2170), .B0 (nx2054), .B1 (
          nx2172)) ;
    xnor2 ix2285 (.Y (nx2284), .A0 (nx2184), .A1 (nx3286)) ;
    oai32 ix2185 (.Y (nx2184), .A0 (nx2643), .A1 (nx1629), .A2 (nx3220), .B0 (
          nx3214), .B1 (nx3216)) ;
    xnor2 ix3287 (.Y (nx3286), .A0 (nx3288), .A1 (nx3290)) ;
    aoi32 ix3289 (.Y (nx3288), .A0 (nx3733), .A1 (nx3699), .A2 (nx2162), .B0 (
          nx2074), .B1 (nx2164)) ;
    xnor2 ix3291 (.Y (nx3290), .A0 (nx3292), .A1 (nx3294)) ;
    nand02 ix3293 (.Y (nx3292), .A0 (nx3729), .A1 (nx3699)) ;
    xnor2 ix3295 (.Y (nx3294), .A0 (nx3296), .A1 (nx3299)) ;
    aoi32 ix3297 (.Y (nx3296), .A0 (nx3737), .A1 (nx3695), .A2 (nx2158), .B0 (
          nx2082), .B1 (nx2160)) ;
    xnor2 ix3300 (.Y (nx3299), .A0 (nx3301), .A1 (nx3303)) ;
    nand02 ix3302 (.Y (nx3301), .A0 (nx3733), .A1 (nx3695)) ;
    xnor2 ix3304 (.Y (nx3303), .A0 (nx2206), .A1 (nx2272)) ;
    oai32 ix2207 (.Y (nx2206), .A0 (nx2193), .A1 (nx1825), .A2 (nx3242), .B0 (
          nx3306), .B1 (nx3238)) ;
    xnor2 ix2273 (.Y (nx2272), .A0 (nx3311), .A1 (nx2270)) ;
    nand02 ix3312 (.Y (nx3311), .A0 (nx3737), .A1 (nx3691)) ;
    xnor2 ix2271 (.Y (nx2270), .A0 (nx3314), .A1 (nx2268)) ;
    aoi32 ix3315 (.Y (nx3314), .A0 (nx3745), .A1 (nx3685), .A2 (nx2150), .B0 (
          nx2098), .B1 (nx2152)) ;
    xnor2 ix2269 (.Y (nx2268), .A0 (nx3317), .A1 (nx2266)) ;
    nand02 ix3318 (.Y (nx3317), .A0 (nx3741), .A1 (nx3687)) ;
    xnor2 ix2267 (.Y (nx2266), .A0 (nx3320), .A1 (nx2264)) ;
    aoi32 ix3321 (.Y (nx3320), .A0 (nx3751), .A1 (nx3681), .A2 (nx2146), .B0 (
          nx2106), .B1 (nx2148)) ;
    xnor2 ix2265 (.Y (nx2264), .A0 (nx3324), .A1 (nx2262)) ;
    nand02 ix3325 (.Y (nx3324), .A0 (nx3745), .A1 (nx3683)) ;
    xnor2 ix2263 (.Y (nx2262), .A0 (nx3327), .A1 (nx2260)) ;
    aoi32 ix3328 (.Y (nx3327), .A0 (nx3755), .A1 (nx3677), .A2 (nx2142), .B0 (
          nx2114), .B1 (nx2144)) ;
    xnor2 ix2261 (.Y (nx2260), .A0 (nx3331), .A1 (nx2258)) ;
    nand02 ix3332 (.Y (nx3331), .A0 (nx3751), .A1 (nx3679)) ;
    xnor2 ix2259 (.Y (nx2258), .A0 (nx3334), .A1 (nx2256)) ;
    aoi32 ix3335 (.Y (nx3334), .A0 (nx3759), .A1 (nx3673), .A2 (nx2138), .B0 (
          nx2122), .B1 (nx2140)) ;
    xnor2 ix2257 (.Y (nx2256), .A0 (nx3338), .A1 (nx2254)) ;
    nand02 ix3339 (.Y (nx3338), .A0 (nx3755), .A1 (nx3673)) ;
    xnor2 ix2255 (.Y (nx2254), .A0 (nx2246), .A1 (nx3346)) ;
    oai32 ix2247 (.Y (nx2246), .A0 (nx2972), .A1 (nx2749), .A2 (nx3278), .B0 (
          nx3342), .B1 (nx3274)) ;
    xnor2 ix3347 (.Y (nx3346), .A0 (nx3348), .A1 (nx3350)) ;
    nand02 ix3349 (.Y (nx3348), .A0 (nx3759), .A1 (nx3669)) ;
    nand02 ix3351 (.Y (nx3350), .A0 (nx3763), .A1 (nx3665)) ;
    xor2 ix2771 (.Y (Product[23]), .A0 (nx2290), .A1 (nx2384)) ;
    oai22 ix2291 (.Y (nx2290), .A0 (nx3281), .A1 (nx3354), .B0 (nx3356), .B1 (
          nx3286)) ;
    inv01 ix3357 (.Y (nx3356), .A (nx2184)) ;
    xnor2 ix2385 (.Y (nx2384), .A0 (nx2296), .A1 (nx3360)) ;
    oai32 ix2297 (.Y (nx2296), .A0 (nx2643), .A1 (nx1605), .A2 (nx3294), .B0 (
          nx3288), .B1 (nx3290)) ;
    xnor2 ix3361 (.Y (nx3360), .A0 (nx2302), .A1 (nx2380)) ;
    oai32 ix2303 (.Y (nx2302), .A0 (nx2479), .A1 (nx1703), .A2 (nx3303), .B0 (
          nx3296), .B1 (nx3299)) ;
    xnor2 ix2381 (.Y (nx2380), .A0 (nx3364), .A1 (nx2378)) ;
    nand02 ix3365 (.Y (nx3364), .A0 (nx3729), .A1 (nx3695)) ;
    xnor2 ix2379 (.Y (nx2378), .A0 (nx3367), .A1 (nx2376)) ;
    aoi32 ix3368 (.Y (nx3367), .A0 (nx3739), .A1 (nx3691), .A2 (nx2270), .B0 (
          nx2206), .B1 (nx2272)) ;
    xnor2 ix2377 (.Y (nx2376), .A0 (nx3370), .A1 (nx2374)) ;
    nand02 ix3371 (.Y (nx3370), .A0 (nx3733), .A1 (nx3691)) ;
    xnor2 ix2375 (.Y (nx2374), .A0 (nx3373), .A1 (nx2372)) ;
    aoi32 ix3374 (.Y (nx3373), .A0 (nx3741), .A1 (nx3687), .A2 (nx2266), .B0 (
          nx2214), .B1 (nx2268)) ;
    xnor2 ix2373 (.Y (nx2372), .A0 (nx3377), .A1 (nx2370)) ;
    nand02 ix3378 (.Y (nx3377), .A0 (nx3739), .A1 (nx3687)) ;
    xnor2 ix2371 (.Y (nx2370), .A0 (nx3380), .A1 (nx2368)) ;
    aoi32 ix3381 (.Y (nx3380), .A0 (nx3747), .A1 (nx3683), .A2 (nx2262), .B0 (
          nx2222), .B1 (nx2264)) ;
    xnor2 ix2369 (.Y (nx2368), .A0 (nx3384), .A1 (nx2366)) ;
    nand02 ix3385 (.Y (nx3384), .A0 (nx3741), .A1 (nx3683)) ;
    xnor2 ix2367 (.Y (nx2366), .A0 (nx3387), .A1 (nx2364)) ;
    aoi32 ix3388 (.Y (nx3387), .A0 (nx3751), .A1 (nx3679), .A2 (nx2258), .B0 (
          nx2230), .B1 (nx2260)) ;
    xnor2 ix2365 (.Y (nx2364), .A0 (nx3391), .A1 (nx2362)) ;
    nand02 ix3392 (.Y (nx3391), .A0 (nx3747), .A1 (nx3679)) ;
    xnor2 ix2363 (.Y (nx2362), .A0 (nx3394), .A1 (nx2360)) ;
    aoi32 ix3395 (.Y (nx3394), .A0 (nx3755), .A1 (nx3673), .A2 (nx2254), .B0 (
          nx2238), .B1 (nx2256)) ;
    xnor2 ix2361 (.Y (nx2360), .A0 (nx3398), .A1 (nx2358)) ;
    nand02 ix3399 (.Y (nx3398), .A0 (nx3751), .A1 (nx3675)) ;
    xnor2 ix2359 (.Y (nx2358), .A0 (nx2350), .A1 (nx3406)) ;
    oai32 ix2351 (.Y (nx2350), .A0 (nx1855), .A1 (nx2749), .A2 (nx3350), .B0 (
          nx3402), .B1 (nx3346)) ;
    xnor2 ix3407 (.Y (nx3406), .A0 (nx3408), .A1 (nx3410)) ;
    nand02 ix3409 (.Y (nx3408), .A0 (nx3755), .A1 (nx3669)) ;
    nand02 ix3411 (.Y (nx3410), .A0 (nx3759), .A1 (nx3665)) ;
    xnor2 ix2769 (.Y (Product[24]), .A0 (nx3413), .A1 (nx2472)) ;
    aoi22 ix3414 (.Y (nx3413), .A0 (nx2296), .A1 (nx2382), .B0 (nx2290), .B1 (
          nx2384)) ;
    xnor2 ix2473 (.Y (nx2472), .A0 (nx3417), .A1 (nx2470)) ;
    aoi32 ix3418 (.Y (nx3417), .A0 (nx3729), .A1 (nx3695), .A2 (nx2378), .B0 (
          nx2302), .B1 (nx2380)) ;
    xnor2 ix2471 (.Y (nx2470), .A0 (nx3420), .A1 (nx2468)) ;
    aoi32 ix3421 (.Y (nx3420), .A0 (nx3733), .A1 (nx3691), .A2 (nx2374), .B0 (
          nx2310), .B1 (nx2376)) ;
    xnor2 ix2469 (.Y (nx2468), .A0 (nx3424), .A1 (nx2466)) ;
    nand02 ix3425 (.Y (nx3424), .A0 (nx3729), .A1 (nx3691)) ;
    xnor2 ix2467 (.Y (nx2466), .A0 (nx3427), .A1 (nx2464)) ;
    aoi32 ix3428 (.Y (nx3427), .A0 (nx3739), .A1 (nx3687), .A2 (nx2370), .B0 (
          nx2318), .B1 (nx2372)) ;
    xnor2 ix2465 (.Y (nx2464), .A0 (nx3431), .A1 (nx2462)) ;
    nand02 ix3432 (.Y (nx3431), .A0 (nx3735), .A1 (nx3687)) ;
    xnor2 ix2463 (.Y (nx2462), .A0 (nx3434), .A1 (nx2460)) ;
    aoi32 ix3435 (.Y (nx3434), .A0 (nx3743), .A1 (nx3683), .A2 (nx2366), .B0 (
          nx2326), .B1 (nx2368)) ;
    xnor2 ix2461 (.Y (nx2460), .A0 (nx3438), .A1 (nx2458)) ;
    nand02 ix3439 (.Y (nx3438), .A0 (nx3739), .A1 (nx3683)) ;
    xnor2 ix2459 (.Y (nx2458), .A0 (nx3441), .A1 (nx2456)) ;
    aoi32 ix3442 (.Y (nx3441), .A0 (nx3747), .A1 (nx3679), .A2 (nx2362), .B0 (
          nx2334), .B1 (nx2364)) ;
    xnor2 ix2457 (.Y (nx2456), .A0 (nx3445), .A1 (nx2454)) ;
    nand02 ix3446 (.Y (nx3445), .A0 (nx3743), .A1 (nx3679)) ;
    xnor2 ix2455 (.Y (nx2454), .A0 (nx3448), .A1 (nx2452)) ;
    aoi32 ix3449 (.Y (nx3448), .A0 (nx3751), .A1 (nx3675), .A2 (nx2358), .B0 (
          nx2342), .B1 (nx2360)) ;
    xnor2 ix2453 (.Y (nx2452), .A0 (nx3452), .A1 (nx2450)) ;
    nand02 ix3453 (.Y (nx3452), .A0 (nx3747), .A1 (nx3675)) ;
    xnor2 ix2451 (.Y (nx2450), .A0 (nx2442), .A1 (nx3460)) ;
    oai32 ix2443 (.Y (nx2442), .A0 (nx1567), .A1 (nx2749), .A2 (nx3410), .B0 (
          nx3456), .B1 (nx3406)) ;
    xnor2 ix3461 (.Y (nx3460), .A0 (nx3462), .A1 (nx3464)) ;
    nand02 ix3463 (.Y (nx3462), .A0 (nx3751), .A1 (nx3669)) ;
    nand02 ix3465 (.Y (nx3464), .A0 (nx3755), .A1 (nx3665)) ;
    xor2 ix2767 (.Y (Product[25]), .A0 (nx2478), .A1 (nx2548)) ;
    oai22 ix2479 (.Y (nx2478), .A0 (nx3413), .A1 (nx3468), .B0 (nx3417), .B1 (
          nx3470)) ;
    xnor2 ix2549 (.Y (nx2548), .A0 (nx3473), .A1 (nx2546)) ;
    aoi32 ix3474 (.Y (nx3473), .A0 (nx3729), .A1 (nx3691), .A2 (nx2466), .B0 (
          nx2402), .B1 (nx2468)) ;
    xnor2 ix2547 (.Y (nx2546), .A0 (nx3477), .A1 (nx2544)) ;
    aoi32 ix3478 (.Y (nx3477), .A0 (nx3735), .A1 (nx3687), .A2 (nx2462), .B0 (
          nx2410), .B1 (nx2464)) ;
    xnor2 ix2545 (.Y (nx2544), .A0 (nx3481), .A1 (nx2542)) ;
    nand02 ix3482 (.Y (nx3481), .A0 (nx3729), .A1 (nx3687)) ;
    xnor2 ix2543 (.Y (nx2542), .A0 (nx3484), .A1 (nx2540)) ;
    aoi32 ix3485 (.Y (nx3484), .A0 (nx3739), .A1 (nx3683), .A2 (nx2458), .B0 (
          nx2418), .B1 (nx2460)) ;
    xnor2 ix2541 (.Y (nx2540), .A0 (nx3488), .A1 (nx2538)) ;
    nand02 ix3489 (.Y (nx3488), .A0 (nx3735), .A1 (nx3683)) ;
    xnor2 ix2539 (.Y (nx2538), .A0 (nx3491), .A1 (nx2536)) ;
    aoi32 ix3492 (.Y (nx3491), .A0 (nx3743), .A1 (nx3679), .A2 (nx2454), .B0 (
          nx2426), .B1 (nx2456)) ;
    xnor2 ix2537 (.Y (nx2536), .A0 (nx3495), .A1 (nx2534)) ;
    nand02 ix3496 (.Y (nx3495), .A0 (nx3739), .A1 (nx3679)) ;
    xnor2 ix2535 (.Y (nx2534), .A0 (nx3498), .A1 (nx2532)) ;
    aoi32 ix3499 (.Y (nx3498), .A0 (nx3747), .A1 (nx3675), .A2 (nx2450), .B0 (
          nx2434), .B1 (nx2452)) ;
    xnor2 ix2533 (.Y (nx2532), .A0 (nx3502), .A1 (nx2530)) ;
    nand02 ix3503 (.Y (nx3502), .A0 (nx3743), .A1 (nx3675)) ;
    xnor2 ix2531 (.Y (nx2530), .A0 (nx2522), .A1 (nx3510)) ;
    oai32 ix2523 (.Y (nx2522), .A0 (nx2948), .A1 (nx2749), .A2 (nx3464), .B0 (
          nx3506), .B1 (nx3460)) ;
    xnor2 ix3511 (.Y (nx3510), .A0 (nx3512), .A1 (nx3514)) ;
    nand02 ix3513 (.Y (nx3512), .A0 (nx3747), .A1 (nx3669)) ;
    nand02 ix3515 (.Y (nx3514), .A0 (nx3751), .A1 (nx3665)) ;
    xnor2 ix2765 (.Y (Product[26]), .A0 (nx3517), .A1 (nx2612)) ;
    aoi22 ix3518 (.Y (nx3517), .A0 (nx2484), .A1 (nx2546), .B0 (nx2478), .B1 (
          nx2548)) ;
    xnor2 ix2613 (.Y (nx2612), .A0 (nx3521), .A1 (nx2610)) ;
    aoi32 ix3522 (.Y (nx3521), .A0 (nx3731), .A1 (nx3687), .A2 (nx2542), .B0 (
          nx2490), .B1 (nx2544)) ;
    xnor2 ix2611 (.Y (nx2610), .A0 (nx3525), .A1 (nx2608)) ;
    aoi32 ix3526 (.Y (nx3525), .A0 (nx3735), .A1 (nx3683), .A2 (nx2538), .B0 (
          nx2498), .B1 (nx2540)) ;
    xnor2 ix2609 (.Y (nx2608), .A0 (nx3529), .A1 (nx2606)) ;
    nand02 ix3530 (.Y (nx3529), .A0 (nx3731), .A1 (nx3683)) ;
    xnor2 ix2607 (.Y (nx2606), .A0 (nx3532), .A1 (nx2604)) ;
    aoi32 ix3533 (.Y (nx3532), .A0 (nx3739), .A1 (nx3679), .A2 (nx2534), .B0 (
          nx2506), .B1 (nx2536)) ;
    xnor2 ix2605 (.Y (nx2604), .A0 (nx3536), .A1 (nx2602)) ;
    nand02 ix3537 (.Y (nx3536), .A0 (nx3735), .A1 (nx3679)) ;
    xnor2 ix2603 (.Y (nx2602), .A0 (nx3539), .A1 (nx2600)) ;
    aoi32 ix3540 (.Y (nx3539), .A0 (nx3743), .A1 (nx3675), .A2 (nx2530), .B0 (
          nx2514), .B1 (nx2532)) ;
    xnor2 ix2601 (.Y (nx2600), .A0 (nx3543), .A1 (nx2598)) ;
    nand02 ix3544 (.Y (nx3543), .A0 (nx3739), .A1 (nx3675)) ;
    xnor2 ix2599 (.Y (nx2598), .A0 (nx2590), .A1 (nx3551)) ;
    oai32 ix2591 (.Y (nx2590), .A0 (nx1559), .A1 (nx2749), .A2 (nx3514), .B0 (
          nx3547), .B1 (nx3510)) ;
    xnor2 ix3552 (.Y (nx3551), .A0 (nx3553), .A1 (nx3555)) ;
    nand02 ix3554 (.Y (nx3553), .A0 (nx3743), .A1 (nx3669)) ;
    nand02 ix3556 (.Y (nx3555), .A0 (nx3747), .A1 (nx3665)) ;
    xor2 ix2763 (.Y (Product[27]), .A0 (nx2618), .A1 (nx2664)) ;
    oai22 ix2619 (.Y (nx2618), .A0 (nx3517), .A1 (nx3559), .B0 (nx3521), .B1 (
          nx3561)) ;
    xnor2 ix2665 (.Y (nx2664), .A0 (nx3564), .A1 (nx2662)) ;
    aoi32 ix3565 (.Y (nx3564), .A0 (nx3731), .A1 (nx3683), .A2 (nx2606), .B0 (
          nx2566), .B1 (nx2608)) ;
    xnor2 ix2663 (.Y (nx2662), .A0 (nx3568), .A1 (nx2660)) ;
    aoi32 ix3569 (.Y (nx3568), .A0 (nx3735), .A1 (nx3679), .A2 (nx2602), .B0 (
          nx2574), .B1 (nx2604)) ;
    xnor2 ix2661 (.Y (nx2660), .A0 (nx3572), .A1 (nx2658)) ;
    nand02 ix3573 (.Y (nx3572), .A0 (nx3731), .A1 (nx3679)) ;
    xnor2 ix2659 (.Y (nx2658), .A0 (nx3575), .A1 (nx2656)) ;
    aoi32 ix3576 (.Y (nx3575), .A0 (nx3739), .A1 (nx3675), .A2 (nx2598), .B0 (
          nx2582), .B1 (nx2600)) ;
    xnor2 ix2657 (.Y (nx2656), .A0 (nx3579), .A1 (nx2654)) ;
    nand02 ix3580 (.Y (nx3579), .A0 (nx3735), .A1 (nx3675)) ;
    xnor2 ix2655 (.Y (nx2654), .A0 (nx2646), .A1 (nx3587)) ;
    oai32 ix2647 (.Y (nx2646), .A0 (nx2193), .A1 (nx2749), .A2 (nx3555), .B0 (
          nx3583), .B1 (nx3551)) ;
    xnor2 ix3588 (.Y (nx3587), .A0 (nx3589), .A1 (nx3591)) ;
    nand02 ix3590 (.Y (nx3589), .A0 (nx3739), .A1 (nx3669)) ;
    nand02 ix3592 (.Y (nx3591), .A0 (nx3743), .A1 (nx3665)) ;
    xnor2 ix2761 (.Y (Product[28]), .A0 (nx3594), .A1 (nx2704)) ;
    aoi22 ix3595 (.Y (nx3594), .A0 (nx2624), .A1 (nx2662), .B0 (nx2618), .B1 (
          nx2664)) ;
    xnor2 ix2705 (.Y (nx2704), .A0 (nx3598), .A1 (nx2702)) ;
    aoi32 ix3599 (.Y (nx3598), .A0 (nx3731), .A1 (nx3679), .A2 (nx2658), .B0 (
          nx2630), .B1 (nx2660)) ;
    xnor2 ix2703 (.Y (nx2702), .A0 (nx3602), .A1 (nx2700)) ;
    aoi32 ix3603 (.Y (nx3602), .A0 (nx3735), .A1 (nx3675), .A2 (nx2654), .B0 (
          nx2638), .B1 (nx2656)) ;
    xnor2 ix2701 (.Y (nx2700), .A0 (nx3606), .A1 (nx2698)) ;
    nand02 ix3607 (.Y (nx3606), .A0 (nx3731), .A1 (nx3675)) ;
    xnor2 ix2699 (.Y (nx2698), .A0 (nx2690), .A1 (nx3614)) ;
    oai32 ix2691 (.Y (nx2690), .A0 (nx2918), .A1 (nx2749), .A2 (nx3591), .B0 (
          nx3610), .B1 (nx3587)) ;
    xnor2 ix3615 (.Y (nx3614), .A0 (nx3616), .A1 (nx3618)) ;
    nand02 ix3617 (.Y (nx3616), .A0 (nx3735), .A1 (nx3671)) ;
    nand02 ix3619 (.Y (nx3618), .A0 (nx3739), .A1 (nx3665)) ;
    xor2 ix2759 (.Y (Product[29]), .A0 (nx2710), .A1 (nx2732)) ;
    oai22 ix2711 (.Y (nx2710), .A0 (nx3594), .A1 (nx3622), .B0 (nx3598), .B1 (
          nx3624)) ;
    xnor2 ix2733 (.Y (nx2732), .A0 (nx3627), .A1 (nx2730)) ;
    aoi32 ix3628 (.Y (nx3627), .A0 (nx3731), .A1 (nx3675), .A2 (nx2698), .B0 (
          nx2682), .B1 (nx2700)) ;
    xnor2 ix2731 (.Y (nx2730), .A0 (nx2722), .A1 (nx3636)) ;
    oai32 ix2723 (.Y (nx2722), .A0 (nx2479), .A1 (nx2749), .A2 (nx3618), .B0 (
          nx3632), .B1 (nx3614)) ;
    xnor2 ix3637 (.Y (nx3636), .A0 (nx3638), .A1 (nx3640)) ;
    nand02 ix3639 (.Y (nx3638), .A0 (nx3731), .A1 (nx3671)) ;
    nand02 ix3641 (.Y (nx3640), .A0 (nx3735), .A1 (nx3667)) ;
    xnor2 ix2751 (.Y (Product[30]), .A0 (nx3643), .A1 (nx2748)) ;
    aoi22 ix3644 (.Y (nx3643), .A0 (nx2716), .A1 (nx2730), .B0 (nx2710), .B1 (
          nx2732)) ;
    xnor2 ix2749 (.Y (nx2748), .A0 (nx2744), .A1 (nx3652)) ;
    oai32 ix2745 (.Y (nx2744), .A0 (nx2643), .A1 (nx2749), .A2 (nx3640), .B0 (
          nx3648), .B1 (nx3636)) ;
    nand02 ix3653 (.Y (nx3652), .A0 (nx3731), .A1 (nx3667)) ;
    ao32 ix2757 (.Y (Product[31]), .A0 (nx2744), .A1 (nx3731), .A2 (nx3667), .B0 (
         nx2738), .B1 (nx2748)) ;
    inv01 ix2739 (.Y (nx2738), .A (nx3643)) ;
    inv01 ix3649 (.Y (nx3648), .A (nx2722)) ;
    inv01 ix2717 (.Y (nx2716), .A (nx3627)) ;
    inv01 ix3623 (.Y (nx3622), .A (nx2704)) ;
    inv01 ix3625 (.Y (nx3624), .A (nx2702)) ;
    inv01 ix3633 (.Y (nx3632), .A (nx2690)) ;
    inv01 ix2683 (.Y (nx2682), .A (nx3602)) ;
    inv01 ix3611 (.Y (nx3610), .A (nx2646)) ;
    inv01 ix2639 (.Y (nx2638), .A (nx3575)) ;
    inv01 ix2631 (.Y (nx2630), .A (nx3568)) ;
    inv01 ix2625 (.Y (nx2624), .A (nx3564)) ;
    inv01 ix3560 (.Y (nx3559), .A (nx2612)) ;
    inv01 ix3562 (.Y (nx3561), .A (nx2610)) ;
    inv01 ix3584 (.Y (nx3583), .A (nx2590)) ;
    inv01 ix2583 (.Y (nx2582), .A (nx3539)) ;
    inv01 ix2575 (.Y (nx2574), .A (nx3532)) ;
    inv01 ix2567 (.Y (nx2566), .A (nx3525)) ;
    inv01 ix3548 (.Y (nx3547), .A (nx2522)) ;
    inv01 ix2515 (.Y (nx2514), .A (nx3498)) ;
    inv01 ix2507 (.Y (nx2506), .A (nx3491)) ;
    inv01 ix2499 (.Y (nx2498), .A (nx3484)) ;
    inv01 ix2491 (.Y (nx2490), .A (nx3477)) ;
    inv01 ix2485 (.Y (nx2484), .A (nx3473)) ;
    inv01 ix3469 (.Y (nx3468), .A (nx2472)) ;
    inv01 ix3471 (.Y (nx3470), .A (nx2470)) ;
    inv01 ix3507 (.Y (nx3506), .A (nx2442)) ;
    inv01 ix2435 (.Y (nx2434), .A (nx3448)) ;
    inv01 ix2427 (.Y (nx2426), .A (nx3441)) ;
    inv01 ix2419 (.Y (nx2418), .A (nx3434)) ;
    inv01 ix2411 (.Y (nx2410), .A (nx3427)) ;
    inv01 ix2403 (.Y (nx2402), .A (nx3420)) ;
    inv01 ix2383 (.Y (nx2382), .A (nx3360)) ;
    inv01 ix3457 (.Y (nx3456), .A (nx2350)) ;
    inv01 ix2343 (.Y (nx2342), .A (nx3394)) ;
    inv01 ix2335 (.Y (nx2334), .A (nx3387)) ;
    inv01 ix2327 (.Y (nx2326), .A (nx3380)) ;
    inv01 ix2319 (.Y (nx2318), .A (nx3373)) ;
    inv01 ix2311 (.Y (nx2310), .A (nx3367)) ;
    inv01 ix3355 (.Y (nx3354), .A (nx2284)) ;
    inv01 ix3403 (.Y (nx3402), .A (nx2246)) ;
    inv01 ix2239 (.Y (nx2238), .A (nx3334)) ;
    inv01 ix2231 (.Y (nx2230), .A (nx3327)) ;
    inv01 ix2223 (.Y (nx2222), .A (nx3320)) ;
    inv01 ix2215 (.Y (nx2214), .A (nx3314)) ;
    inv01 ix2171 (.Y (nx2170), .A (nx3212)) ;
    inv01 ix3343 (.Y (nx3342), .A (nx2130)) ;
    inv01 ix2123 (.Y (nx2122), .A (nx3262)) ;
    inv01 ix2115 (.Y (nx2114), .A (nx3255)) ;
    inv01 ix2107 (.Y (nx2106), .A (nx3249)) ;
    inv01 ix3307 (.Y (nx3306), .A (nx2090)) ;
    inv01 ix2083 (.Y (nx2082), .A (nx3229)) ;
    inv01 ix3205 (.Y (nx3204), .A (nx2048)) ;
    inv01 ix3271 (.Y (nx3270), .A (nx2002)) ;
    inv01 ix1995 (.Y (nx1994), .A (nx3184)) ;
    inv01 ix1987 (.Y (nx1986), .A (nx3178)) ;
    inv01 ix3207 (.Y (nx3206), .A (nx1924)) ;
    inv01 ix3193 (.Y (nx3192), .A (nx1862)) ;
    inv01 ix1855 (.Y (nx1854), .A (nx3102)) ;
    inv01 ix3124 (.Y (nx3123), .A (nx1782)) ;
    inv01 ix1777 (.Y (nx1776), .A (nx3028)) ;
    inv01 ix3024 (.Y (nx3023), .A (nx1764)) ;
    inv01 ix3026 (.Y (nx3025), .A (nx1762)) ;
    inv01 ix3110 (.Y (nx3109), .A (nx1710)) ;
    inv01 ix3083 (.Y (nx3082), .A (nx1678)) ;
    inv01 ix1671 (.Y (nx1670), .A (nx2964)) ;
    inv01 ix1663 (.Y (nx1662), .A (nx2958)) ;
    inv01 ix3034 (.Y (nx3033), .A (nx1630)) ;
    inv01 ix1623 (.Y (nx1622), .A (nx2910)) ;
    inv01 ix1603 (.Y (nx1602), .A (nx2787)) ;
    inv01 ix3005 (.Y (nx3004), .A (nx1546)) ;
    inv01 ix1539 (.Y (nx1538), .A (nx2875)) ;
    inv01 ix2975 (.Y (nx2974), .A (nx1522)) ;
    inv01 ix1515 (.Y (nx1514), .A (nx2849)) ;
    inv01 ix2951 (.Y (nx2950), .A (nx1498)) ;
    inv01 ix1491 (.Y (nx1490), .A (nx2823)) ;
    inv01 ix2921 (.Y (nx2920), .A (nx1474)) ;
    inv01 ix1467 (.Y (nx1466), .A (nx2797)) ;
    inv01 ix1447 (.Y (nx1446), .A (nx2775)) ;
    inv01 ix1441 (.Y (nx1440), .A (nx2639)) ;
    inv01 ix1383 (.Y (nx1382), .A (nx3007)) ;
    inv01 ix2884 (.Y (nx2883), .A (nx1370)) ;
    inv01 ix1263 (.Y (nx1262), .A (nx2637)) ;
    inv01 ix2746 (.Y (nx2745), .A (nx1196)) ;
    inv01 ix2576 (.Y (nx2575), .A (nx1032)) ;
    inv01 ix2388 (.Y (nx2387), .A (nx880)) ;
    inv01 ix2162 (.Y (nx2161), .A (nx740)) ;
    inv01 ix1976 (.Y (nx1975), .A (nx612)) ;
    inv01 ix1822 (.Y (nx1821), .A (nx496)) ;
    inv01 ix1700 (.Y (nx1699), .A (nx392)) ;
    inv01 ix1602 (.Y (nx1601), .A (nx300)) ;
    inv01 ix1662 (.Y (nx1661), .A (nx220)) ;
    inv01 ix1758 (.Y (nx1757), .A (nx152)) ;
    inv01 ix1888 (.Y (nx1887), .A (nx96)) ;
    inv01 ix2048 (.Y (nx2047), .A (nx52)) ;
    inv01 ix2248 (.Y (nx2247), .A (nx20)) ;
    and02 ix3 (.Y (Product[0]), .A0 (nx3791), .A1 (nx3727)) ;
    inv01 ix3664 (.Y (nx3665), .A (nx2761)) ;
    inv01 ix3666 (.Y (nx3667), .A (nx2761)) ;
    inv01 ix3668 (.Y (nx3669), .A (nx2749)) ;
    inv01 ix3670 (.Y (nx3671), .A (nx2749)) ;
    inv01 ix3672 (.Y (nx3673), .A (nx2579)) ;
    inv01 ix3674 (.Y (nx3675), .A (nx2579)) ;
    inv01 ix3676 (.Y (nx3677), .A (nx2391)) ;
    inv01 ix3678 (.Y (nx3679), .A (nx2391)) ;
    inv01 ix3680 (.Y (nx3681), .A (nx2165)) ;
    inv01 ix3682 (.Y (nx3683), .A (nx2165)) ;
    inv01 ix3684 (.Y (nx3685), .A (nx1979)) ;
    inv01 ix3686 (.Y (nx3687), .A (nx1979)) ;
    inv01 ix3688 (.Y (nx3689), .A (nx1825)) ;
    inv01 ix3690 (.Y (nx3691), .A (nx1825)) ;
    inv01 ix3692 (.Y (nx3693), .A (nx1703)) ;
    inv01 ix3694 (.Y (nx3695), .A (nx1703)) ;
    inv01 ix3696 (.Y (nx3697), .A (nx1605)) ;
    inv01 ix3698 (.Y (nx3699), .A (nx1605)) ;
    inv01 ix3700 (.Y (nx3701), .A (nx1629)) ;
    inv01 ix3702 (.Y (nx3703), .A (nx1629)) ;
    inv01 ix3704 (.Y (nx3705), .A (nx1589)) ;
    inv01 ix3706 (.Y (nx3707), .A (nx1589)) ;
    inv01 ix3708 (.Y (nx3709), .A (nx1581)) ;
    inv01 ix3710 (.Y (nx3711), .A (nx1581)) ;
    inv01 ix3712 (.Y (nx3713), .A (nx1733)) ;
    inv01 ix3714 (.Y (nx3715), .A (nx1733)) ;
    inv01 ix3716 (.Y (nx3717), .A (nx1569)) ;
    inv01 ix3718 (.Y (nx3719), .A (nx1569)) ;
    inv01 ix3720 (.Y (nx3721), .A (nx1561)) ;
    inv01 ix3722 (.Y (nx3723), .A (nx1561)) ;
    inv01 ix3724 (.Y (nx3725), .A (nx2195)) ;
    inv01 ix3726 (.Y (nx3727), .A (nx2195)) ;
    inv01 ix3728 (.Y (nx3729), .A (nx2643)) ;
    inv01 ix3730 (.Y (nx3731), .A (nx2643)) ;
    inv01 ix3732 (.Y (nx3733), .A (nx2479)) ;
    inv01 ix3734 (.Y (nx3735), .A (nx2479)) ;
    inv01 ix3736 (.Y (nx3737), .A (nx2918)) ;
    inv01 ix3738 (.Y (nx3739), .A (nx2918)) ;
    inv01 ix3740 (.Y (nx3741), .A (nx2193)) ;
    inv01 ix3742 (.Y (nx3743), .A (nx2193)) ;
    inv01 ix3744 (.Y (nx3745), .A (nx1559)) ;
    inv01 ix3746 (.Y (nx3747), .A (nx1559)) ;
    inv01 ix3748 (.Y (nx3749), .A (nx2948)) ;
    inv01 ix3750 (.Y (nx3751), .A (nx2948)) ;
    inv01 ix3752 (.Y (nx3753), .A (nx1567)) ;
    inv01 ix3754 (.Y (nx3755), .A (nx1567)) ;
    inv01 ix3756 (.Y (nx3757), .A (nx1855)) ;
    inv01 ix3758 (.Y (nx3759), .A (nx1855)) ;
    inv01 ix3760 (.Y (nx3761), .A (nx2972)) ;
    inv01 ix3762 (.Y (nx3763), .A (nx2972)) ;
    inv01 ix3764 (.Y (nx3765), .A (nx1731)) ;
    inv01 ix3766 (.Y (nx3767), .A (nx1731)) ;
    inv01 ix3768 (.Y (nx3769), .A (nx1579)) ;
    inv01 ix3770 (.Y (nx3771), .A (nx1579)) ;
    inv01 ix3772 (.Y (nx3773), .A (nx3002)) ;
    inv01 ix3774 (.Y (nx3775), .A (nx3002)) ;
    inv01 ix3776 (.Y (nx3777), .A (nx1587)) ;
    inv01 ix3778 (.Y (nx3779), .A (nx1587)) ;
    inv01 ix3780 (.Y (nx3781), .A (nx1627)) ;
    inv01 ix3782 (.Y (nx3783), .A (nx1627)) ;
    inv01 ix3784 (.Y (nx3785), .A (nx1631)) ;
    inv01 ix3786 (.Y (nx3787), .A (nx1631)) ;
    inv01 ix3788 (.Y (nx3789), .A (nx1607)) ;
    inv01 ix3790 (.Y (nx3791), .A (nx1607)) ;
endmodule

